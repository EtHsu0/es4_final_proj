library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity eight_segments is
    port (
        row : in unsigned (9 downto 0);
        col : in unsigned (9 downto 0);
        clk : in std_logic;
        rgb : out std_logic_vector(5 downto 0)
    );
end eight_segments;

architecture synth of eight_segments is
    signal addr : std_logic_vector(13 downto 0);

    begin
        addr <= std_logic_vector(row(7 downto 0)) & std_logic_vector(col(7 downto 0));
        process(clk) is begin
            if rising_edge(clk) then 
                case addr is 
                when "00000000000000" => rgb <= "000000";
                when "00000000000001" => rgb <= "000000";
                when "00000000000010" => rgb <= "000000";
                when "00000000000011" => rgb <= "000000";
                when "00000000000100" => rgb <= "000000";
                when "00000000000101" => rgb <= "000000";
                when "00000000000110" => rgb <= "000000";
                when "00000000000111" => rgb <= "000000";
                when "00000000001000" => rgb <= "000000";
                when "00000000001001" => rgb <= "000000";
                when "00000000001010" => rgb <= "000000";
                when "00000000001011" => rgb <= "000000";
                when "00000000001100" => rgb <= "000000";
                when "00000000001101" => rgb <= "000000";
                when "00000000001110" => rgb <= "000000";
                when "00000000001111" => rgb <= "000000";
                when "00000000010000" => rgb <= "000000";
                when "00000000010001" => rgb <= "000000";
                when "00000000010010" => rgb <= "000000";
                when "00000000010011" => rgb <= "000000";
                when "00000000010100" => rgb <= "000000";
                when "00000000010101" => rgb <= "000000";
                when "00000000010110" => rgb <= "000000";
                when "00000000010111" => rgb <= "000000";
                when "00000000011000" => rgb <= "000000";
                when "00000000011001" => rgb <= "000000";
                when "00000000011010" => rgb <= "010000";
                when "00000000011011" => rgb <= "010000";
                when "00000000011100" => rgb <= "010000";
                when "00000000011101" => rgb <= "000000";
                when "00000000011110" => rgb <= "000000";
                when "00000000011111" => rgb <= "000000";
                when "00000000100000" => rgb <= "000000";
                when "00000000100001" => rgb <= "000000";
                when "00000000100010" => rgb <= "000000";
                when "00000000100011" => rgb <= "000000";
                when "00000000100100" => rgb <= "000000";
                when "00000000100101" => rgb <= "000000";
                when "00000000100110" => rgb <= "000000";
                when "00000000100111" => rgb <= "000000";
                when "00000000101000" => rgb <= "000000";
                when "00000000101001" => rgb <= "000000";
                when "00000000101010" => rgb <= "000000";
                when "00000000101011" => rgb <= "000000";
                when "00000010000000" => rgb <= "000000";
                when "00000010000001" => rgb <= "000000";
                when "00000010000010" => rgb <= "000000";
                when "00000010000011" => rgb <= "000000";
                when "00000010000100" => rgb <= "000000";
                when "00000010000101" => rgb <= "000000";
                when "00000010000110" => rgb <= "000000";
                when "00000010000111" => rgb <= "000000";
                when "00000010001000" => rgb <= "000000";
                when "00000010001001" => rgb <= "000000";
                when "00000010001010" => rgb <= "000000";
                when "00000010001011" => rgb <= "000000";
                when "00000010001100" => rgb <= "000000";
                when "00000010001101" => rgb <= "000000";
                when "00000010001110" => rgb <= "000000";
                when "00000010001111" => rgb <= "000000";
                when "00000010010000" => rgb <= "000000";
                when "00000010010001" => rgb <= "000000";
                when "00000010010010" => rgb <= "000000";
                when "00000010010011" => rgb <= "000000";
                when "00000010010100" => rgb <= "000000";
                when "00000010010101" => rgb <= "000000";
                when "00000010010110" => rgb <= "000000";
                when "00000010010111" => rgb <= "000000";
                when "00000010011000" => rgb <= "000000";
                when "00000010011001" => rgb <= "000000";
                when "00000010011010" => rgb <= "010000";
                when "00000010011011" => rgb <= "010000";
                when "00000010011100" => rgb <= "010000";
                when "00000010011101" => rgb <= "000000";
                when "00000010011110" => rgb <= "000000";
                when "00000010011111" => rgb <= "000000";
                when "00000010100000" => rgb <= "000000";
                when "00000010100001" => rgb <= "000000";
                when "00000010100010" => rgb <= "000000";
                when "00000010100011" => rgb <= "000000";
                when "00000010100100" => rgb <= "000000";
                when "00000010100101" => rgb <= "000000";
                when "00000010100110" => rgb <= "000000";
                when "00000010100111" => rgb <= "000000";
                when "00000010101000" => rgb <= "000000";
                when "00000010101001" => rgb <= "000000";
                when "00000010101010" => rgb <= "000000";
                when "00000010101011" => rgb <= "000000";
                when "00000100000000" => rgb <= "000000";
                when "00000100000001" => rgb <= "000000";
                when "00000100000010" => rgb <= "000000";
                when "00000100000011" => rgb <= "000000";
                when "00000100000100" => rgb <= "000000";
                when "00000100000101" => rgb <= "000000";
                when "00000100000110" => rgb <= "000000";
                when "00000100000111" => rgb <= "000000";
                when "00000100001000" => rgb <= "000000";
                when "00000100001001" => rgb <= "000000";
                when "00000100001010" => rgb <= "000000";
                when "00000100001011" => rgb <= "000000";
                when "00000100001100" => rgb <= "000000";
                when "00000100001101" => rgb <= "000000";
                when "00000100001110" => rgb <= "000000";
                when "00000100001111" => rgb <= "000000";
                when "00000100010000" => rgb <= "000000";
                when "00000100010001" => rgb <= "000000";
                when "00000100010010" => rgb <= "000000";
                when "00000100010011" => rgb <= "000000";
                when "00000100010100" => rgb <= "000000";
                when "00000100010101" => rgb <= "000000";
                when "00000100010110" => rgb <= "000000";
                when "00000100010111" => rgb <= "000000";
                when "00000100011000" => rgb <= "000000";
                when "00000100011001" => rgb <= "000000";
                when "00000100011010" => rgb <= "010000";
                when "00000100011011" => rgb <= "010000";
                when "00000100011100" => rgb <= "010000";
                when "00000100011101" => rgb <= "000000";
                when "00000100011110" => rgb <= "000000";
                when "00000100011111" => rgb <= "000000";
                when "00000100100000" => rgb <= "000000";
                when "00000100100001" => rgb <= "000000";
                when "00000100100010" => rgb <= "000000";
                when "00000100100011" => rgb <= "000000";
                when "00000100100100" => rgb <= "000000";
                when "00000100100101" => rgb <= "000000";
                when "00000100100110" => rgb <= "000000";
                when "00000100100111" => rgb <= "000000";
                when "00000100101000" => rgb <= "000000";
                when "00000100101001" => rgb <= "000000";
                when "00000100101010" => rgb <= "000000";
                when "00000100101011" => rgb <= "000000";
                when "00000110000000" => rgb <= "000000";
                when "00000110000001" => rgb <= "000000";
                when "00000110000010" => rgb <= "000000";
                when "00000110000011" => rgb <= "000000";
                when "00000110000100" => rgb <= "000000";
                when "00000110000101" => rgb <= "000000";
                when "00000110000110" => rgb <= "000000";
                when "00000110000111" => rgb <= "000000";
                when "00000110001000" => rgb <= "000000";
                when "00000110001001" => rgb <= "000000";
                when "00000110001010" => rgb <= "000000";
                when "00000110001011" => rgb <= "000000";
                when "00000110001100" => rgb <= "000000";
                when "00000110001101" => rgb <= "000000";
                when "00000110001110" => rgb <= "000000";
                when "00000110001111" => rgb <= "000000";
                when "00000110010000" => rgb <= "000000";
                when "00000110010001" => rgb <= "000000";
                when "00000110010010" => rgb <= "000000";
                when "00000110010011" => rgb <= "000000";
                when "00000110010100" => rgb <= "000000";
                when "00000110010101" => rgb <= "000000";
                when "00000110010110" => rgb <= "010000";
                when "00000110010111" => rgb <= "010000";
                when "00000110011000" => rgb <= "010000";
                when "00000110011001" => rgb <= "010000";
                when "00000110011010" => rgb <= "010000";
                when "00000110011011" => rgb <= "010000";
                when "00000110011100" => rgb <= "010000";
                when "00000110011101" => rgb <= "000000";
                when "00000110011110" => rgb <= "000000";
                when "00000110011111" => rgb <= "000000";
                when "00000110100000" => rgb <= "000000";
                when "00000110100001" => rgb <= "000000";
                when "00000110100010" => rgb <= "000000";
                when "00000110100011" => rgb <= "000000";
                when "00000110100100" => rgb <= "000000";
                when "00000110100101" => rgb <= "000000";
                when "00000110100110" => rgb <= "000000";
                when "00000110100111" => rgb <= "000000";
                when "00000110101000" => rgb <= "000000";
                when "00000110101001" => rgb <= "000000";
                when "00000110101010" => rgb <= "000000";
                when "00000110101011" => rgb <= "000000";
                when "00001000000000" => rgb <= "000000";
                when "00001000000001" => rgb <= "000000";
                when "00001000000010" => rgb <= "000000";
                when "00001000000011" => rgb <= "000000";
                when "00001000000100" => rgb <= "000000";
                when "00001000000101" => rgb <= "000000";
                when "00001000000110" => rgb <= "000000";
                when "00001000000111" => rgb <= "000000";
                when "00001000001000" => rgb <= "000000";
                when "00001000001001" => rgb <= "000000";
                when "00001000001010" => rgb <= "000000";
                when "00001000001011" => rgb <= "000000";
                when "00001000001100" => rgb <= "000000";
                when "00001000001101" => rgb <= "000000";
                when "00001000001110" => rgb <= "000000";
                when "00001000001111" => rgb <= "000000";
                when "00001000010000" => rgb <= "000000";
                when "00001000010001" => rgb <= "000000";
                when "00001000010010" => rgb <= "000000";
                when "00001000010011" => rgb <= "000000";
                when "00001000010100" => rgb <= "000000";
                when "00001000010101" => rgb <= "000000";
                when "00001000010110" => rgb <= "010000";
                when "00001000010111" => rgb <= "010000";
                when "00001000011000" => rgb <= "010000";
                when "00001000011001" => rgb <= "010000";
                when "00001000011010" => rgb <= "000000";
                when "00001000011011" => rgb <= "000000";
                when "00001000011100" => rgb <= "000000";
                when "00001000011101" => rgb <= "000000";
                when "00001000011110" => rgb <= "000000";
                when "00001000011111" => rgb <= "000000";
                when "00001000100000" => rgb <= "000000";
                when "00001000100001" => rgb <= "000000";
                when "00001000100010" => rgb <= "000000";
                when "00001000100011" => rgb <= "000000";
                when "00001000100100" => rgb <= "000000";
                when "00001000100101" => rgb <= "000000";
                when "00001000100110" => rgb <= "000000";
                when "00001000100111" => rgb <= "000000";
                when "00001000101000" => rgb <= "000000";
                when "00001000101001" => rgb <= "000000";
                when "00001000101010" => rgb <= "000000";
                when "00001000101011" => rgb <= "000000";
                when "00001010000000" => rgb <= "000000";
                when "00001010000001" => rgb <= "000000";
                when "00001010000010" => rgb <= "000000";
                when "00001010000011" => rgb <= "000000";
                when "00001010000100" => rgb <= "000000";
                when "00001010000101" => rgb <= "000000";
                when "00001010000110" => rgb <= "000000";
                when "00001010000111" => rgb <= "000000";
                when "00001010001000" => rgb <= "000000";
                when "00001010001001" => rgb <= "000000";
                when "00001010001010" => rgb <= "000000";
                when "00001010001011" => rgb <= "000000";
                when "00001010001100" => rgb <= "000000";
                when "00001010001101" => rgb <= "000000";
                when "00001010001110" => rgb <= "000000";
                when "00001010001111" => rgb <= "000000";
                when "00001010010000" => rgb <= "000000";
                when "00001010010001" => rgb <= "000000";
                when "00001010010010" => rgb <= "000000";
                when "00001010010011" => rgb <= "000000";
                when "00001010010100" => rgb <= "000000";
                when "00001010010101" => rgb <= "000000";
                when "00001010010110" => rgb <= "010000";
                when "00001010010111" => rgb <= "010000";
                when "00001010011000" => rgb <= "010000";
                when "00001010011001" => rgb <= "010000";
                when "00001010011010" => rgb <= "000000";
                when "00001010011011" => rgb <= "000000";
                when "00001010011100" => rgb <= "000000";
                when "00001010011101" => rgb <= "000000";
                when "00001010011110" => rgb <= "000000";
                when "00001010011111" => rgb <= "000000";
                when "00001010100000" => rgb <= "000000";
                when "00001010100001" => rgb <= "000000";
                when "00001010100010" => rgb <= "000000";
                when "00001010100011" => rgb <= "000000";
                when "00001010100100" => rgb <= "000000";
                when "00001010100101" => rgb <= "000000";
                when "00001010100110" => rgb <= "000000";
                when "00001010100111" => rgb <= "000000";
                when "00001010101000" => rgb <= "000000";
                when "00001010101001" => rgb <= "000000";
                when "00001010101010" => rgb <= "000000";
                when "00001010101011" => rgb <= "000000";
                when "00001100000000" => rgb <= "000000";
                when "00001100000001" => rgb <= "000000";
                when "00001100000010" => rgb <= "000000";
                when "00001100000011" => rgb <= "000000";
                when "00001100000100" => rgb <= "000000";
                when "00001100000101" => rgb <= "000000";
                when "00001100000110" => rgb <= "000000";
                when "00001100000111" => rgb <= "000000";
                when "00001100001000" => rgb <= "000000";
                when "00001100001001" => rgb <= "000000";
                when "00001100001010" => rgb <= "000000";
                when "00001100001011" => rgb <= "100101";
                when "00001100001100" => rgb <= "100101";
                when "00001100001101" => rgb <= "100101";
                when "00001100001110" => rgb <= "100101";
                when "00001100001111" => rgb <= "100100";
                when "00001100010000" => rgb <= "100100";
                when "00001100010001" => rgb <= "100100";
                when "00001100010010" => rgb <= "010000";
                when "00001100010011" => rgb <= "010000";
                when "00001100010100" => rgb <= "010000";
                when "00001100010101" => rgb <= "010000";
                when "00001100010110" => rgb <= "010000";
                when "00001100010111" => rgb <= "010000";
                when "00001100011000" => rgb <= "010000";
                when "00001100011001" => rgb <= "010000";
                when "00001100011010" => rgb <= "010000";
                when "00001100011011" => rgb <= "010000";
                when "00001100011100" => rgb <= "010001";
                when "00001100011101" => rgb <= "010001";
                when "00001100011110" => rgb <= "010001";
                when "00001100011111" => rgb <= "010001";
                when "00001100100000" => rgb <= "010001";
                when "00001100100001" => rgb <= "000000";
                when "00001100100010" => rgb <= "000000";
                when "00001100100011" => rgb <= "000000";
                when "00001100100100" => rgb <= "000000";
                when "00001100100101" => rgb <= "000000";
                when "00001100100110" => rgb <= "000000";
                when "00001100100111" => rgb <= "000000";
                when "00001100101000" => rgb <= "000000";
                when "00001100101001" => rgb <= "000000";
                when "00001100101010" => rgb <= "000000";
                when "00001100101011" => rgb <= "000000";
                when "00001110000000" => rgb <= "000000";
                when "00001110000001" => rgb <= "000000";
                when "00001110000010" => rgb <= "000000";
                when "00001110000011" => rgb <= "000000";
                when "00001110000100" => rgb <= "000000";
                when "00001110000101" => rgb <= "000000";
                when "00001110000110" => rgb <= "000000";
                when "00001110000111" => rgb <= "000000";
                when "00001110001000" => rgb <= "000000";
                when "00001110001001" => rgb <= "000000";
                when "00001110001010" => rgb <= "000000";
                when "00001110001011" => rgb <= "100101";
                when "00001110001100" => rgb <= "100101";
                when "00001110001101" => rgb <= "100101";
                when "00001110001110" => rgb <= "100100";
                when "00001110001111" => rgb <= "100100";
                when "00001110010000" => rgb <= "100100";
                when "00001110010001" => rgb <= "100100";
                when "00001110010010" => rgb <= "010000";
                when "00001110010011" => rgb <= "010000";
                when "00001110010100" => rgb <= "010000";
                when "00001110010101" => rgb <= "010000";
                when "00001110010110" => rgb <= "010000";
                when "00001110010111" => rgb <= "010000";
                when "00001110011000" => rgb <= "010000";
                when "00001110011001" => rgb <= "010000";
                when "00001110011010" => rgb <= "010001";
                when "00001110011011" => rgb <= "010001";
                when "00001110011100" => rgb <= "010001";
                when "00001110011101" => rgb <= "010001";
                when "00001110011110" => rgb <= "010001";
                when "00001110011111" => rgb <= "010001";
                when "00001110100000" => rgb <= "010001";
                when "00001110100001" => rgb <= "000000";
                when "00001110100010" => rgb <= "000000";
                when "00001110100011" => rgb <= "000000";
                when "00001110100100" => rgb <= "000000";
                when "00001110100101" => rgb <= "000000";
                when "00001110100110" => rgb <= "000000";
                when "00001110100111" => rgb <= "000000";
                when "00001110101000" => rgb <= "000000";
                when "00001110101001" => rgb <= "000000";
                when "00001110101010" => rgb <= "000000";
                when "00001110101011" => rgb <= "000000";
                when "00010000000000" => rgb <= "000000";
                when "00010000000001" => rgb <= "000000";
                when "00010000000010" => rgb <= "000000";
                when "00010000000011" => rgb <= "000000";
                when "00010000000100" => rgb <= "000000";
                when "00010000000101" => rgb <= "000000";
                when "00010000000110" => rgb <= "000000";
                when "00010000000111" => rgb <= "000000";
                when "00010000001000" => rgb <= "000000";
                when "00010000001001" => rgb <= "000000";
                when "00010000001010" => rgb <= "000000";
                when "00010000001011" => rgb <= "100101";
                when "00010000001100" => rgb <= "100101";
                when "00010000001101" => rgb <= "100101";
                when "00010000001110" => rgb <= "100101";
                when "00010000001111" => rgb <= "100100";
                when "00010000010000" => rgb <= "100100";
                when "00010000010001" => rgb <= "100100";
                when "00010000010010" => rgb <= "010000";
                when "00010000010011" => rgb <= "010000";
                when "00010000010100" => rgb <= "010000";
                when "00010000010101" => rgb <= "010000";
                when "00010000010110" => rgb <= "010000";
                when "00010000010111" => rgb <= "010000";
                when "00010000011000" => rgb <= "010001";
                when "00010000011001" => rgb <= "010001";
                when "00010000011010" => rgb <= "010001";
                when "00010000011011" => rgb <= "010001";
                when "00010000011100" => rgb <= "010001";
                when "00010000011101" => rgb <= "010001";
                when "00010000011110" => rgb <= "010001";
                when "00010000011111" => rgb <= "010001";
                when "00010000100000" => rgb <= "010001";
                when "00010000100001" => rgb <= "000000";
                when "00010000100010" => rgb <= "000000";
                when "00010000100011" => rgb <= "000000";
                when "00010000100100" => rgb <= "000000";
                when "00010000100101" => rgb <= "000000";
                when "00010000100110" => rgb <= "000000";
                when "00010000100111" => rgb <= "000000";
                when "00010000101000" => rgb <= "000000";
                when "00010000101001" => rgb <= "000000";
                when "00010000101010" => rgb <= "000000";
                when "00010000101011" => rgb <= "000000";
                when "00010010000000" => rgb <= "000000";
                when "00010010000001" => rgb <= "000000";
                when "00010010000010" => rgb <= "000000";
                when "00010010000011" => rgb <= "000000";
                when "00010010000100" => rgb <= "000000";
                when "00010010000101" => rgb <= "000000";
                when "00010010000110" => rgb <= "000000";
                when "00010010000111" => rgb <= "000000";
                when "00010010001000" => rgb <= "000000";
                when "00010010001001" => rgb <= "000000";
                when "00010010001010" => rgb <= "000000";
                when "00010010001011" => rgb <= "101001";
                when "00010010001100" => rgb <= "100101";
                when "00010010001101" => rgb <= "100101";
                when "00010010001110" => rgb <= "100101";
                when "00010010001111" => rgb <= "100100";
                when "00010010010000" => rgb <= "100100";
                when "00010010010001" => rgb <= "100100";
                when "00010010010010" => rgb <= "010000";
                when "00010010010011" => rgb <= "010000";
                when "00010010010100" => rgb <= "010000";
                when "00010010010101" => rgb <= "010000";
                when "00010010010110" => rgb <= "010000";
                when "00010010010111" => rgb <= "010001";
                when "00010010011000" => rgb <= "010001";
                when "00010010011001" => rgb <= "010101";
                when "00010010011010" => rgb <= "100101";
                when "00010010011011" => rgb <= "100101";
                when "00010010011100" => rgb <= "100101";
                when "00010010011101" => rgb <= "100101";
                when "00010010011110" => rgb <= "100101";
                when "00010010011111" => rgb <= "100101";
                when "00010010100000" => rgb <= "100101";
                when "00010010100001" => rgb <= "000000";
                when "00010010100010" => rgb <= "000000";
                when "00010010100011" => rgb <= "000000";
                when "00010010100100" => rgb <= "000000";
                when "00010010100101" => rgb <= "000000";
                when "00010010100110" => rgb <= "000000";
                when "00010010100111" => rgb <= "000000";
                when "00010010101000" => rgb <= "000000";
                when "00010010101001" => rgb <= "000000";
                when "00010010101010" => rgb <= "000000";
                when "00010010101011" => rgb <= "000000";
                when "00010100000000" => rgb <= "000000";
                when "00010100000001" => rgb <= "000000";
                when "00010100000010" => rgb <= "000000";
                when "00010100000011" => rgb <= "000000";
                when "00010100000100" => rgb <= "100101";
                when "00010100000101" => rgb <= "100101";
                when "00010100000110" => rgb <= "100101";
                when "00010100000111" => rgb <= "100101";
                when "00010100001000" => rgb <= "101001";
                when "00010100001001" => rgb <= "101001";
                when "00010100001010" => rgb <= "101001";
                when "00010100001011" => rgb <= "111010";
                when "00010100001100" => rgb <= "111010";
                when "00010100001101" => rgb <= "111010";
                when "00010100001110" => rgb <= "101010";
                when "00010100001111" => rgb <= "101001";
                when "00010100010000" => rgb <= "101000";
                when "00010100010001" => rgb <= "101000";
                when "00010100010010" => rgb <= "010000";
                when "00010100010011" => rgb <= "010000";
                when "00010100010100" => rgb <= "010000";
                when "00010100010101" => rgb <= "010000";
                when "00010100010110" => rgb <= "100101";
                when "00010100010111" => rgb <= "100101";
                when "00010100011000" => rgb <= "100101";
                when "00010100011001" => rgb <= "100101";
                when "00010100011010" => rgb <= "111010";
                when "00010100011011" => rgb <= "111010";
                when "00010100011100" => rgb <= "111010";
                when "00010100011101" => rgb <= "101001";
                when "00010100011110" => rgb <= "111001";
                when "00010100011111" => rgb <= "111001";
                when "00010100100000" => rgb <= "111001";
                when "00010100100001" => rgb <= "010001";
                when "00010100100010" => rgb <= "010001";
                when "00010100100011" => rgb <= "010001";
                when "00010100100100" => rgb <= "010001";
                when "00010100100101" => rgb <= "010001";
                when "00010100100110" => rgb <= "010001";
                when "00010100100111" => rgb <= "010001";
                when "00010100101000" => rgb <= "000000";
                when "00010100101001" => rgb <= "000000";
                when "00010100101010" => rgb <= "000000";
                when "00010100101011" => rgb <= "000000";
                when "00010110000000" => rgb <= "000000";
                when "00010110000001" => rgb <= "000000";
                when "00010110000010" => rgb <= "000000";
                when "00010110000011" => rgb <= "000000";
                when "00010110000100" => rgb <= "100101";
                when "00010110000101" => rgb <= "100101";
                when "00010110000110" => rgb <= "100101";
                when "00010110000111" => rgb <= "100101";
                when "00010110001000" => rgb <= "101001";
                when "00010110001001" => rgb <= "101001";
                when "00010110001010" => rgb <= "101001";
                when "00010110001011" => rgb <= "111010";
                when "00010110001100" => rgb <= "111111";
                when "00010110001101" => rgb <= "111111";
                when "00010110001110" => rgb <= "101010";
                when "00010110001111" => rgb <= "101001";
                when "00010110010000" => rgb <= "101001";
                when "00010110010001" => rgb <= "101001";
                when "00010110010010" => rgb <= "010000";
                when "00010110010011" => rgb <= "010000";
                when "00010110010100" => rgb <= "010000";
                when "00010110010101" => rgb <= "010000";
                when "00010110010110" => rgb <= "100101";
                when "00010110010111" => rgb <= "100101";
                when "00010110011000" => rgb <= "100101";
                when "00010110011001" => rgb <= "100101";
                when "00010110011010" => rgb <= "111010";
                when "00010110011011" => rgb <= "111010";
                when "00010110011100" => rgb <= "111010";
                when "00010110011101" => rgb <= "101001";
                when "00010110011110" => rgb <= "111001";
                when "00010110011111" => rgb <= "111001";
                when "00010110100000" => rgb <= "111001";
                when "00010110100001" => rgb <= "010001";
                when "00010110100010" => rgb <= "010001";
                when "00010110100011" => rgb <= "010001";
                when "00010110100100" => rgb <= "010001";
                when "00010110100101" => rgb <= "010001";
                when "00010110100110" => rgb <= "010001";
                when "00010110100111" => rgb <= "010001";
                when "00010110101000" => rgb <= "000000";
                when "00010110101001" => rgb <= "000000";
                when "00010110101010" => rgb <= "000000";
                when "00010110101011" => rgb <= "000000";
                when "00011000000000" => rgb <= "000000";
                when "00011000000001" => rgb <= "000000";
                when "00011000000010" => rgb <= "000000";
                when "00011000000011" => rgb <= "000000";
                when "00011000000100" => rgb <= "100101";
                when "00011000000101" => rgb <= "100101";
                when "00011000000110" => rgb <= "100101";
                when "00011000000111" => rgb <= "100101";
                when "00011000001000" => rgb <= "101001";
                when "00011000001001" => rgb <= "101001";
                when "00011000001010" => rgb <= "101001";
                when "00011000001011" => rgb <= "111010";
                when "00011000001100" => rgb <= "111110";
                when "00011000001101" => rgb <= "111110";
                when "00011000001110" => rgb <= "101010";
                when "00011000001111" => rgb <= "101001";
                when "00011000010000" => rgb <= "101001";
                when "00011000010001" => rgb <= "101001";
                when "00011000010010" => rgb <= "010000";
                when "00011000010011" => rgb <= "010000";
                when "00011000010100" => rgb <= "010000";
                when "00011000010101" => rgb <= "010000";
                when "00011000010110" => rgb <= "100101";
                when "00011000010111" => rgb <= "100101";
                when "00011000011000" => rgb <= "100101";
                when "00011000011001" => rgb <= "100101";
                when "00011000011010" => rgb <= "101010";
                when "00011000011011" => rgb <= "101010";
                when "00011000011100" => rgb <= "101010";
                when "00011000011101" => rgb <= "101001";
                when "00011000011110" => rgb <= "101001";
                when "00011000011111" => rgb <= "101001";
                when "00011000100000" => rgb <= "101001";
                when "00011000100001" => rgb <= "010001";
                when "00011000100010" => rgb <= "010001";
                when "00011000100011" => rgb <= "010001";
                when "00011000100100" => rgb <= "010001";
                when "00011000100101" => rgb <= "010001";
                when "00011000100110" => rgb <= "010001";
                when "00011000100111" => rgb <= "010001";
                when "00011000101000" => rgb <= "000000";
                when "00011000101001" => rgb <= "000000";
                when "00011000101010" => rgb <= "000000";
                when "00011000101011" => rgb <= "000000";
                when "00011010000000" => rgb <= "100101";
                when "00011010000001" => rgb <= "100101";
                when "00011010000010" => rgb <= "100101";
                when "00011010000011" => rgb <= "100101";
                when "00011010000100" => rgb <= "100101";
                when "00011010000101" => rgb <= "100101";
                when "00011010000110" => rgb <= "100101";
                when "00011010000111" => rgb <= "101001";
                when "00011010001000" => rgb <= "101001";
                when "00011010001001" => rgb <= "101001";
                when "00011010001010" => rgb <= "101001";
                when "00011010001011" => rgb <= "101010";
                when "00011010001100" => rgb <= "101110";
                when "00011010001101" => rgb <= "101110";
                when "00011010001110" => rgb <= "101010";
                when "00011010001111" => rgb <= "101010";
                when "00011010010000" => rgb <= "101010";
                when "00011010010001" => rgb <= "101010";
                when "00011010010010" => rgb <= "101010";
                when "00011010010011" => rgb <= "101010";
                when "00011010010100" => rgb <= "101010";
                when "00011010010101" => rgb <= "101010";
                when "00011010010110" => rgb <= "101010";
                when "00011010010111" => rgb <= "101010";
                when "00011010011000" => rgb <= "101010";
                when "00011010011001" => rgb <= "101010";
                when "00011010011010" => rgb <= "111010";
                when "00011010011011" => rgb <= "111010";
                when "00011010011100" => rgb <= "111010";
                when "00011010011101" => rgb <= "101010";
                when "00011010011110" => rgb <= "101010";
                when "00011010011111" => rgb <= "101010";
                when "00011010100000" => rgb <= "101010";
                when "00011010100001" => rgb <= "100101";
                when "00011010100010" => rgb <= "100101";
                when "00011010100011" => rgb <= "100101";
                when "00011010100100" => rgb <= "100101";
                when "00011010100101" => rgb <= "010001";
                when "00011010100110" => rgb <= "010001";
                when "00011010100111" => rgb <= "010001";
                when "00011010101000" => rgb <= "010001";
                when "00011010101001" => rgb <= "010001";
                when "00011010101010" => rgb <= "010001";
                when "00011010101011" => rgb <= "010001";
                when "00011100000000" => rgb <= "100101";
                when "00011100000001" => rgb <= "100101";
                when "00011100000010" => rgb <= "100101";
                when "00011100000011" => rgb <= "100101";
                when "00011100000100" => rgb <= "101001";
                when "00011100000101" => rgb <= "101001";
                when "00011100000110" => rgb <= "101001";
                when "00011100000111" => rgb <= "101001";
                when "00011100001000" => rgb <= "101001";
                when "00011100001001" => rgb <= "101001";
                when "00011100001010" => rgb <= "101010";
                when "00011100001011" => rgb <= "111110";
                when "00011100001100" => rgb <= "101110";
                when "00011100001101" => rgb <= "101110";
                when "00011100001110" => rgb <= "101010";
                when "00011100001111" => rgb <= "111010";
                when "00011100010000" => rgb <= "111111";
                when "00011100010001" => rgb <= "101110";
                when "00011100010010" => rgb <= "101110";
                when "00011100010011" => rgb <= "101110";
                when "00011100010100" => rgb <= "101010";
                when "00011100010101" => rgb <= "111010";
                when "00011100010110" => rgb <= "101011";
                when "00011100010111" => rgb <= "111011";
                when "00011100011000" => rgb <= "111011";
                when "00011100011001" => rgb <= "101110";
                when "00011100011010" => rgb <= "111110";
                when "00011100011011" => rgb <= "111110";
                when "00011100011100" => rgb <= "111110";
                when "00011100011101" => rgb <= "101010";
                when "00011100011110" => rgb <= "101010";
                when "00011100011111" => rgb <= "111010";
                when "00011100100000" => rgb <= "111010";
                when "00011100100001" => rgb <= "101001";
                when "00011100100010" => rgb <= "101001";
                when "00011100100011" => rgb <= "101001";
                when "00011100100100" => rgb <= "100101";
                when "00011100100101" => rgb <= "010001";
                when "00011100100110" => rgb <= "010001";
                when "00011100100111" => rgb <= "010001";
                when "00011100101000" => rgb <= "010001";
                when "00011100101001" => rgb <= "010001";
                when "00011100101010" => rgb <= "010001";
                when "00011100101011" => rgb <= "010001";
                when "00011110000000" => rgb <= "100101";
                when "00011110000001" => rgb <= "100101";
                when "00011110000010" => rgb <= "100101";
                when "00011110000011" => rgb <= "100101";
                when "00011110000100" => rgb <= "101001";
                when "00011110000101" => rgb <= "101001";
                when "00011110000110" => rgb <= "101001";
                when "00011110000111" => rgb <= "101001";
                when "00011110001000" => rgb <= "101001";
                when "00011110001001" => rgb <= "101001";
                when "00011110001010" => rgb <= "101010";
                when "00011110001011" => rgb <= "111110";
                when "00011110001100" => rgb <= "111110";
                when "00011110001101" => rgb <= "111010";
                when "00011110001110" => rgb <= "101110";
                when "00011110001111" => rgb <= "111110";
                when "00011110010000" => rgb <= "111110";
                when "00011110010001" => rgb <= "101110";
                when "00011110010010" => rgb <= "111111";
                when "00011110010011" => rgb <= "111110";
                when "00011110010100" => rgb <= "101110";
                when "00011110010101" => rgb <= "111011";
                when "00011110010110" => rgb <= "101010";
                when "00011110010111" => rgb <= "111010";
                when "00011110011000" => rgb <= "111010";
                when "00011110011001" => rgb <= "111110";
                when "00011110011010" => rgb <= "111110";
                when "00011110011011" => rgb <= "111110";
                when "00011110011100" => rgb <= "111010";
                when "00011110011101" => rgb <= "101010";
                when "00011110011110" => rgb <= "101010";
                when "00011110011111" => rgb <= "101010";
                when "00011110100000" => rgb <= "101010";
                when "00011110100001" => rgb <= "101001";
                when "00011110100010" => rgb <= "101001";
                when "00011110100011" => rgb <= "101001";
                when "00011110100100" => rgb <= "100101";
                when "00011110100101" => rgb <= "010001";
                when "00011110100110" => rgb <= "010001";
                when "00011110100111" => rgb <= "010001";
                when "00011110101000" => rgb <= "010000";
                when "00011110101001" => rgb <= "010000";
                when "00011110101010" => rgb <= "010000";
                when "00011110101011" => rgb <= "010000";
                when "00100000000000" => rgb <= "100101";
                when "00100000000001" => rgb <= "100101";
                when "00100000000010" => rgb <= "100101";
                when "00100000000011" => rgb <= "100101";
                when "00100000000100" => rgb <= "101001";
                when "00100000000101" => rgb <= "101001";
                when "00100000000110" => rgb <= "101001";
                when "00100000000111" => rgb <= "101001";
                when "00100000001000" => rgb <= "101010";
                when "00100000001001" => rgb <= "101010";
                when "00100000001010" => rgb <= "101010";
                when "00100000001011" => rgb <= "111010";
                when "00100000001100" => rgb <= "111010";
                when "00100000001101" => rgb <= "111010";
                when "00100000001110" => rgb <= "111010";
                when "00100000001111" => rgb <= "111010";
                when "00100000010000" => rgb <= "111010";
                when "00100000010001" => rgb <= "111010";
                when "00100000010010" => rgb <= "111010";
                when "00100000010011" => rgb <= "111010";
                when "00100000010100" => rgb <= "111010";
                when "00100000010101" => rgb <= "111110";
                when "00100000010110" => rgb <= "111110";
                when "00100000010111" => rgb <= "101110";
                when "00100000011000" => rgb <= "101110";
                when "00100000011001" => rgb <= "101110";
                when "00100000011010" => rgb <= "101110";
                when "00100000011011" => rgb <= "101110";
                when "00100000011100" => rgb <= "101110";
                when "00100000011101" => rgb <= "101010";
                when "00100000011110" => rgb <= "111010";
                when "00100000011111" => rgb <= "111010";
                when "00100000100000" => rgb <= "111001";
                when "00100000100001" => rgb <= "101001";
                when "00100000100010" => rgb <= "101001";
                when "00100000100011" => rgb <= "101001";
                when "00100000100100" => rgb <= "100101";
                when "00100000100101" => rgb <= "010000";
                when "00100000100110" => rgb <= "010000";
                when "00100000100111" => rgb <= "010000";
                when "00100000101000" => rgb <= "010000";
                when "00100000101001" => rgb <= "010000";
                when "00100000101010" => rgb <= "010000";
                when "00100000101011" => rgb <= "010000";
                when "00100010000000" => rgb <= "100101";
                when "00100010000001" => rgb <= "100101";
                when "00100010000010" => rgb <= "100101";
                when "00100010000011" => rgb <= "100101";
                when "00100010000100" => rgb <= "101001";
                when "00100010000101" => rgb <= "101001";
                when "00100010000110" => rgb <= "101001";
                when "00100010000111" => rgb <= "101001";
                when "00100010001000" => rgb <= "101010";
                when "00100010001001" => rgb <= "111010";
                when "00100010001010" => rgb <= "101010";
                when "00100010001011" => rgb <= "101110";
                when "00100010001100" => rgb <= "101110";
                when "00100010001101" => rgb <= "101010";
                when "00100010001110" => rgb <= "111010";
                when "00100010001111" => rgb <= "111010";
                when "00100010010000" => rgb <= "101010";
                when "00100010010001" => rgb <= "101010";
                when "00100010010010" => rgb <= "101010";
                when "00100010010011" => rgb <= "101010";
                when "00100010010100" => rgb <= "101010";
                when "00100010010101" => rgb <= "101010";
                when "00100010010110" => rgb <= "101010";
                when "00100010010111" => rgb <= "101010";
                when "00100010011000" => rgb <= "101010";
                when "00100010011001" => rgb <= "101010";
                when "00100010011010" => rgb <= "101010";
                when "00100010011011" => rgb <= "101010";
                when "00100010011100" => rgb <= "101010";
                when "00100010011101" => rgb <= "101001";
                when "00100010011110" => rgb <= "101001";
                when "00100010011111" => rgb <= "101001";
                when "00100010100000" => rgb <= "101001";
                when "00100010100001" => rgb <= "101001";
                when "00100010100010" => rgb <= "101001";
                when "00100010100011" => rgb <= "101001";
                when "00100010100100" => rgb <= "101001";
                when "00100010100101" => rgb <= "101001";
                when "00100010100110" => rgb <= "101001";
                when "00100010100111" => rgb <= "101001";
                when "00100010101000" => rgb <= "100101";
                when "00100010101001" => rgb <= "010000";
                when "00100010101010" => rgb <= "010000";
                when "00100010101011" => rgb <= "010000";
                when "00100100000000" => rgb <= "100101";
                when "00100100000001" => rgb <= "100101";
                when "00100100000010" => rgb <= "100101";
                when "00100100000011" => rgb <= "100101";
                when "00100100000100" => rgb <= "101001";
                when "00100100000101" => rgb <= "101001";
                when "00100100000110" => rgb <= "101001";
                when "00100100000111" => rgb <= "101001";
                when "00100100001000" => rgb <= "111010";
                when "00100100001001" => rgb <= "101010";
                when "00100100001010" => rgb <= "101010";
                when "00100100001011" => rgb <= "101010";
                when "00100100001100" => rgb <= "101010";
                when "00100100001101" => rgb <= "111110";
                when "00100100001110" => rgb <= "111110";
                when "00100100001111" => rgb <= "111110";
                when "00100100010000" => rgb <= "111010";
                when "00100100010001" => rgb <= "111110";
                when "00100100010010" => rgb <= "101110";
                when "00100100010011" => rgb <= "101110";
                when "00100100010100" => rgb <= "111110";
                when "00100100010101" => rgb <= "111010";
                when "00100100010110" => rgb <= "111010";
                when "00100100010111" => rgb <= "111010";
                when "00100100011000" => rgb <= "111010";
                when "00100100011001" => rgb <= "111010";
                when "00100100011010" => rgb <= "101010";
                when "00100100011011" => rgb <= "101001";
                when "00100100011100" => rgb <= "101001";
                when "00100100011101" => rgb <= "101001";
                when "00100100011110" => rgb <= "111001";
                when "00100100011111" => rgb <= "111001";
                when "00100100100000" => rgb <= "101001";
                when "00100100100001" => rgb <= "101001";
                when "00100100100010" => rgb <= "101001";
                when "00100100100011" => rgb <= "111001";
                when "00100100100100" => rgb <= "101001";
                when "00100100100101" => rgb <= "101001";
                when "00100100100110" => rgb <= "101001";
                when "00100100100111" => rgb <= "101001";
                when "00100100101000" => rgb <= "100100";
                when "00100100101001" => rgb <= "010000";
                when "00100100101010" => rgb <= "010000";
                when "00100100101011" => rgb <= "010000";
                when "00100110000000" => rgb <= "100101";
                when "00100110000001" => rgb <= "100101";
                when "00100110000010" => rgb <= "100101";
                when "00100110000011" => rgb <= "100101";
                when "00100110000100" => rgb <= "101001";
                when "00100110000101" => rgb <= "101001";
                when "00100110000110" => rgb <= "101001";
                when "00100110000111" => rgb <= "101001";
                when "00100110001000" => rgb <= "101010";
                when "00100110001001" => rgb <= "101010";
                when "00100110001010" => rgb <= "111010";
                when "00100110001011" => rgb <= "111010";
                when "00100110001100" => rgb <= "111010";
                when "00100110001101" => rgb <= "111010";
                when "00100110001110" => rgb <= "111110";
                when "00100110001111" => rgb <= "111110";
                when "00100110010000" => rgb <= "101110";
                when "00100110010001" => rgb <= "101110";
                when "00100110010010" => rgb <= "101110";
                when "00100110010011" => rgb <= "111010";
                when "00100110010100" => rgb <= "111010";
                when "00100110010101" => rgb <= "101010";
                when "00100110010110" => rgb <= "101010";
                when "00100110010111" => rgb <= "101010";
                when "00100110011000" => rgb <= "101010";
                when "00100110011001" => rgb <= "111010";
                when "00100110011010" => rgb <= "101001";
                when "00100110011011" => rgb <= "101001";
                when "00100110011100" => rgb <= "101001";
                when "00100110011101" => rgb <= "101001";
                when "00100110011110" => rgb <= "111001";
                when "00100110011111" => rgb <= "101001";
                when "00100110100000" => rgb <= "101001";
                when "00100110100001" => rgb <= "111001";
                when "00100110100010" => rgb <= "101001";
                when "00100110100011" => rgb <= "101001";
                when "00100110100100" => rgb <= "101001";
                when "00100110100101" => rgb <= "101001";
                when "00100110100110" => rgb <= "101001";
                when "00100110100111" => rgb <= "101001";
                when "00100110101000" => rgb <= "100100";
                when "00100110101001" => rgb <= "010000";
                when "00100110101010" => rgb <= "010000";
                when "00100110101011" => rgb <= "010000";
                when "00101000000000" => rgb <= "100101";
                when "00101000000001" => rgb <= "100101";
                when "00101000000010" => rgb <= "100101";
                when "00101000000011" => rgb <= "100101";
                when "00101000000100" => rgb <= "101001";
                when "00101000000101" => rgb <= "101001";
                when "00101000000110" => rgb <= "101001";
                when "00101000000111" => rgb <= "101001";
                when "00101000001000" => rgb <= "101010";
                when "00101000001001" => rgb <= "101010";
                when "00101000001010" => rgb <= "101010";
                when "00101000001011" => rgb <= "101010";
                when "00101000001100" => rgb <= "111010";
                when "00101000001101" => rgb <= "111010";
                when "00101000001110" => rgb <= "101010";
                when "00101000001111" => rgb <= "101010";
                when "00101000010000" => rgb <= "101010";
                when "00101000010001" => rgb <= "101010";
                when "00101000010010" => rgb <= "101010";
                when "00101000010011" => rgb <= "111010";
                when "00101000010100" => rgb <= "101010";
                when "00101000010101" => rgb <= "111010";
                when "00101000010110" => rgb <= "101001";
                when "00101000010111" => rgb <= "101001";
                when "00101000011000" => rgb <= "111001";
                when "00101000011001" => rgb <= "111001";
                when "00101000011010" => rgb <= "101001";
                when "00101000011011" => rgb <= "101001";
                when "00101000011100" => rgb <= "101001";
                when "00101000011101" => rgb <= "101001";
                when "00101000011110" => rgb <= "111001";
                when "00101000011111" => rgb <= "111001";
                when "00101000100000" => rgb <= "101001";
                when "00101000100001" => rgb <= "111001";
                when "00101000100010" => rgb <= "101001";
                when "00101000100011" => rgb <= "101001";
                when "00101000100100" => rgb <= "101001";
                when "00101000100101" => rgb <= "101001";
                when "00101000100110" => rgb <= "101001";
                when "00101000100111" => rgb <= "101001";
                when "00101000101000" => rgb <= "010101";
                when "00101000101001" => rgb <= "010000";
                when "00101000101010" => rgb <= "010000";
                when "00101000101011" => rgb <= "010000";
                when "00101010000000" => rgb <= "100101";
                when "00101010000001" => rgb <= "100101";
                when "00101010000010" => rgb <= "100101";
                when "00101010000011" => rgb <= "100101";
                when "00101010000100" => rgb <= "101001";
                when "00101010000101" => rgb <= "101001";
                when "00101010000110" => rgb <= "101001";
                when "00101010000111" => rgb <= "101001";
                when "00101010001000" => rgb <= "111010";
                when "00101010001001" => rgb <= "101010";
                when "00101010001010" => rgb <= "101010";
                when "00101010001011" => rgb <= "101010";
                when "00101010001100" => rgb <= "111010";
                when "00101010001101" => rgb <= "111010";
                when "00101010001110" => rgb <= "101010";
                when "00101010001111" => rgb <= "101010";
                when "00101010010000" => rgb <= "101010";
                when "00101010010001" => rgb <= "101010";
                when "00101010010010" => rgb <= "101010";
                when "00101010010011" => rgb <= "101010";
                when "00101010010100" => rgb <= "101010";
                when "00101010010101" => rgb <= "111010";
                when "00101010010110" => rgb <= "101001";
                when "00101010010111" => rgb <= "101001";
                when "00101010011000" => rgb <= "111001";
                when "00101010011001" => rgb <= "111001";
                when "00101010011010" => rgb <= "111001";
                when "00101010011011" => rgb <= "111001";
                when "00101010011100" => rgb <= "111001";
                when "00101010011101" => rgb <= "111001";
                when "00101010011110" => rgb <= "111001";
                when "00101010011111" => rgb <= "101001";
                when "00101010100000" => rgb <= "101001";
                when "00101010100001" => rgb <= "111001";
                when "00101010100010" => rgb <= "101001";
                when "00101010100011" => rgb <= "101001";
                when "00101010100100" => rgb <= "101001";
                when "00101010100101" => rgb <= "101001";
                when "00101010100110" => rgb <= "101001";
                when "00101010100111" => rgb <= "111001";
                when "00101010101000" => rgb <= "010001";
                when "00101010101001" => rgb <= "010000";
                when "00101010101010" => rgb <= "010000";
                when "00101010101011" => rgb <= "010000";
                when "00101100000000" => rgb <= "100101";
                when "00101100000001" => rgb <= "100101";
                when "00101100000010" => rgb <= "100101";
                when "00101100000011" => rgb <= "100101";
                when "00101100000100" => rgb <= "101001";
                when "00101100000101" => rgb <= "101001";
                when "00101100000110" => rgb <= "101001";
                when "00101100000111" => rgb <= "101010";
                when "00101100001000" => rgb <= "111010";
                when "00101100001001" => rgb <= "111010";
                when "00101100001010" => rgb <= "101010";
                when "00101100001011" => rgb <= "111010";
                when "00101100001100" => rgb <= "111010";
                when "00101100001101" => rgb <= "111010";
                when "00101100001110" => rgb <= "101010";
                when "00101100001111" => rgb <= "101010";
                when "00101100010000" => rgb <= "101010";
                when "00101100010001" => rgb <= "101010";
                when "00101100010010" => rgb <= "101010";
                when "00101100010011" => rgb <= "101010";
                when "00101100010100" => rgb <= "101010";
                when "00101100010101" => rgb <= "111010";
                when "00101100010110" => rgb <= "101001";
                when "00101100010111" => rgb <= "111001";
                when "00101100011000" => rgb <= "111001";
                when "00101100011001" => rgb <= "111001";
                when "00101100011010" => rgb <= "111001";
                when "00101100011011" => rgb <= "111001";
                when "00101100011100" => rgb <= "111001";
                when "00101100011101" => rgb <= "111001";
                when "00101100011110" => rgb <= "111001";
                when "00101100011111" => rgb <= "101001";
                when "00101100100000" => rgb <= "101001";
                when "00101100100001" => rgb <= "111001";
                when "00101100100010" => rgb <= "101001";
                when "00101100100011" => rgb <= "111001";
                when "00101100100100" => rgb <= "101001";
                when "00101100100101" => rgb <= "101001";
                when "00101100100110" => rgb <= "101001";
                when "00101100100111" => rgb <= "111001";
                when "00101100101000" => rgb <= "010001";
                when "00101100101001" => rgb <= "010000";
                when "00101100101010" => rgb <= "010000";
                when "00101100101011" => rgb <= "010000";
                when "00101110000000" => rgb <= "100101";
                when "00101110000001" => rgb <= "100101";
                when "00101110000010" => rgb <= "100101";
                when "00101110000011" => rgb <= "100101";
                when "00101110000100" => rgb <= "111001";
                when "00101110000101" => rgb <= "111001";
                when "00101110000110" => rgb <= "101001";
                when "00101110000111" => rgb <= "101010";
                when "00101110001000" => rgb <= "101010";
                when "00101110001001" => rgb <= "111010";
                when "00101110001010" => rgb <= "101010";
                when "00101110001011" => rgb <= "111010";
                when "00101110001100" => rgb <= "111010";
                when "00101110001101" => rgb <= "111010";
                when "00101110001110" => rgb <= "101010";
                when "00101110001111" => rgb <= "101010";
                when "00101110010000" => rgb <= "111010";
                when "00101110010001" => rgb <= "101010";
                when "00101110010010" => rgb <= "111010";
                when "00101110010011" => rgb <= "101010";
                when "00101110010100" => rgb <= "101001";
                when "00101110010101" => rgb <= "111001";
                when "00101110010110" => rgb <= "101001";
                when "00101110010111" => rgb <= "111001";
                when "00101110011000" => rgb <= "101001";
                when "00101110011001" => rgb <= "101001";
                when "00101110011010" => rgb <= "101001";
                when "00101110011011" => rgb <= "101001";
                when "00101110011100" => rgb <= "101001";
                when "00101110011101" => rgb <= "111001";
                when "00101110011110" => rgb <= "111001";
                when "00101110011111" => rgb <= "111001";
                when "00101110100000" => rgb <= "101001";
                when "00101110100001" => rgb <= "111001";
                when "00101110100010" => rgb <= "101001";
                when "00101110100011" => rgb <= "111001";
                when "00101110100100" => rgb <= "101001";
                when "00101110100101" => rgb <= "101001";
                when "00101110100110" => rgb <= "101001";
                when "00101110100111" => rgb <= "101001";
                when "00101110101000" => rgb <= "010001";
                when "00101110101001" => rgb <= "010000";
                when "00101110101010" => rgb <= "010000";
                when "00101110101011" => rgb <= "010000";
                when "00110000000000" => rgb <= "010001";
                when "00110000000001" => rgb <= "010001";
                when "00110000000010" => rgb <= "010001";
                when "00110000000011" => rgb <= "100101";
                when "00110000000100" => rgb <= "111001";
                when "00110000000101" => rgb <= "101001";
                when "00110000000110" => rgb <= "101001";
                when "00110000000111" => rgb <= "101001";
                when "00110000001000" => rgb <= "101001";
                when "00110000001001" => rgb <= "101001";
                when "00110000001010" => rgb <= "101001";
                when "00110000001011" => rgb <= "101010";
                when "00110000001100" => rgb <= "101010";
                when "00110000001101" => rgb <= "101010";
                when "00110000001110" => rgb <= "101010";
                when "00110000001111" => rgb <= "111010";
                when "00110000010000" => rgb <= "111010";
                when "00110000010001" => rgb <= "101010";
                when "00110000010010" => rgb <= "101001";
                when "00110000010011" => rgb <= "101001";
                when "00110000010100" => rgb <= "101001";
                when "00110000010101" => rgb <= "101001";
                when "00110000010110" => rgb <= "101001";
                when "00110000010111" => rgb <= "101001";
                when "00110000011000" => rgb <= "101000";
                when "00110000011001" => rgb <= "101001";
                when "00110000011010" => rgb <= "111001";
                when "00110000011011" => rgb <= "111001";
                when "00110000011100" => rgb <= "111001";
                when "00110000011101" => rgb <= "101001";
                when "00110000011110" => rgb <= "101000";
                when "00110000011111" => rgb <= "101000";
                when "00110000100000" => rgb <= "101000";
                when "00110000100001" => rgb <= "111001";
                when "00110000100010" => rgb <= "111001";
                when "00110000100011" => rgb <= "111001";
                when "00110000100100" => rgb <= "101001";
                when "00110000100101" => rgb <= "101001";
                when "00110000100110" => rgb <= "101001";
                when "00110000100111" => rgb <= "111001";
                when "00110000101000" => rgb <= "010001";
                when "00110000101001" => rgb <= "010000";
                when "00110000101010" => rgb <= "010000";
                when "00110000101011" => rgb <= "010000";
                when "00110010000000" => rgb <= "010001";
                when "00110010000001" => rgb <= "010001";
                when "00110010000010" => rgb <= "010001";
                when "00110010000011" => rgb <= "100101";
                when "00110010000100" => rgb <= "111001";
                when "00110010000101" => rgb <= "101001";
                when "00110010000110" => rgb <= "101001";
                when "00110010000111" => rgb <= "101001";
                when "00110010001000" => rgb <= "101001";
                when "00110010001001" => rgb <= "111001";
                when "00110010001010" => rgb <= "101001";
                when "00110010001011" => rgb <= "111010";
                when "00110010001100" => rgb <= "111010";
                when "00110010001101" => rgb <= "111010";
                when "00110010001110" => rgb <= "111010";
                when "00110010001111" => rgb <= "111010";
                when "00110010010000" => rgb <= "101010";
                when "00110010010001" => rgb <= "101010";
                when "00110010010010" => rgb <= "101001";
                when "00110010010011" => rgb <= "101001";
                when "00110010010100" => rgb <= "101001";
                when "00110010010101" => rgb <= "101001";
                when "00110010010110" => rgb <= "101000";
                when "00110010010111" => rgb <= "101000";
                when "00110010011000" => rgb <= "101000";
                when "00110010011001" => rgb <= "101001";
                when "00110010011010" => rgb <= "101001";
                when "00110010011011" => rgb <= "111001";
                when "00110010011100" => rgb <= "111001";
                when "00110010011101" => rgb <= "101001";
                when "00110010011110" => rgb <= "101000";
                when "00110010011111" => rgb <= "101000";
                when "00110010100000" => rgb <= "101000";
                when "00110010100001" => rgb <= "111001";
                when "00110010100010" => rgb <= "111001";
                when "00110010100011" => rgb <= "111001";
                when "00110010100100" => rgb <= "101001";
                when "00110010100101" => rgb <= "101001";
                when "00110010100110" => rgb <= "101001";
                when "00110010100111" => rgb <= "111001";
                when "00110010101000" => rgb <= "010001";
                when "00110010101001" => rgb <= "010000";
                when "00110010101010" => rgb <= "010000";
                when "00110010101011" => rgb <= "010000";
                when "00110100000000" => rgb <= "010001";
                when "00110100000001" => rgb <= "010001";
                when "00110100000010" => rgb <= "010001";
                when "00110100000011" => rgb <= "100101";
                when "00110100000100" => rgb <= "101001";
                when "00110100000101" => rgb <= "101001";
                when "00110100000110" => rgb <= "101001";
                when "00110100000111" => rgb <= "101001";
                when "00110100001000" => rgb <= "101001";
                when "00110100001001" => rgb <= "101001";
                when "00110100001010" => rgb <= "101001";
                when "00110100001011" => rgb <= "111010";
                when "00110100001100" => rgb <= "111010";
                when "00110100001101" => rgb <= "111010";
                when "00110100001110" => rgb <= "111010";
                when "00110100001111" => rgb <= "111010";
                when "00110100010000" => rgb <= "101010";
                when "00110100010001" => rgb <= "101001";
                when "00110100010010" => rgb <= "101001";
                when "00110100010011" => rgb <= "101001";
                when "00110100010100" => rgb <= "101001";
                when "00110100010101" => rgb <= "101001";
                when "00110100010110" => rgb <= "101000";
                when "00110100010111" => rgb <= "101000";
                when "00110100011000" => rgb <= "101000";
                when "00110100011001" => rgb <= "101001";
                when "00110100011010" => rgb <= "101001";
                when "00110100011011" => rgb <= "101001";
                when "00110100011100" => rgb <= "101001";
                when "00110100011101" => rgb <= "101001";
                when "00110100011110" => rgb <= "101000";
                when "00110100011111" => rgb <= "101000";
                when "00110100100000" => rgb <= "101000";
                when "00110100100001" => rgb <= "111001";
                when "00110100100010" => rgb <= "111001";
                when "00110100100011" => rgb <= "111001";
                when "00110100100100" => rgb <= "101001";
                when "00110100100101" => rgb <= "101001";
                when "00110100100110" => rgb <= "101001";
                when "00110100100111" => rgb <= "101001";
                when "00110100101000" => rgb <= "010001";
                when "00110100101001" => rgb <= "010000";
                when "00110100101010" => rgb <= "010000";
                when "00110100101011" => rgb <= "010000";
                when "00110110000000" => rgb <= "100001";
                when "00110110000001" => rgb <= "100001";
                when "00110110000010" => rgb <= "100001";
                when "00110110000011" => rgb <= "100101";
                when "00110110000100" => rgb <= "111010";
                when "00110110000101" => rgb <= "101001";
                when "00110110000110" => rgb <= "111001";
                when "00110110000111" => rgb <= "101001";
                when "00110110001000" => rgb <= "101001";
                when "00110110001001" => rgb <= "111001";
                when "00110110001010" => rgb <= "101001";
                when "00110110001011" => rgb <= "101010";
                when "00110110001100" => rgb <= "101010";
                when "00110110001101" => rgb <= "101010";
                when "00110110001110" => rgb <= "101010";
                when "00110110001111" => rgb <= "101010";
                when "00110110010000" => rgb <= "101001";
                when "00110110010001" => rgb <= "101001";
                when "00110110010010" => rgb <= "101001";
                when "00110110010011" => rgb <= "101001";
                when "00110110010100" => rgb <= "101001";
                when "00110110010101" => rgb <= "101000";
                when "00110110010110" => rgb <= "101001";
                when "00110110010111" => rgb <= "101000";
                when "00110110011000" => rgb <= "101000";
                when "00110110011001" => rgb <= "101001";
                when "00110110011010" => rgb <= "101001";
                when "00110110011011" => rgb <= "101001";
                when "00110110011100" => rgb <= "101001";
                when "00110110011101" => rgb <= "101001";
                when "00110110011110" => rgb <= "101000";
                when "00110110011111" => rgb <= "101000";
                when "00110110100000" => rgb <= "101000";
                when "00110110100001" => rgb <= "111001";
                when "00110110100010" => rgb <= "111001";
                when "00110110100011" => rgb <= "111001";
                when "00110110100100" => rgb <= "101001";
                when "00110110100101" => rgb <= "101001";
                when "00110110100110" => rgb <= "101001";
                when "00110110100111" => rgb <= "101001";
                when "00110110101000" => rgb <= "010001";
                when "00110110101001" => rgb <= "010000";
                when "00110110101010" => rgb <= "010000";
                when "00110110101011" => rgb <= "010000";
                when "00111000000000" => rgb <= "100001";
                when "00111000000001" => rgb <= "100001";
                when "00111000000010" => rgb <= "100001";
                when "00111000000011" => rgb <= "100101";
                when "00111000000100" => rgb <= "111010";
                when "00111000000101" => rgb <= "101001";
                when "00111000000110" => rgb <= "111001";
                when "00111000000111" => rgb <= "111001";
                when "00111000001000" => rgb <= "111001";
                when "00111000001001" => rgb <= "111001";
                when "00111000001010" => rgb <= "111001";
                when "00111000001011" => rgb <= "101001";
                when "00111000001100" => rgb <= "101001";
                when "00111000001101" => rgb <= "101001";
                when "00111000001110" => rgb <= "101001";
                when "00111000001111" => rgb <= "101001";
                when "00111000010000" => rgb <= "101001";
                when "00111000010001" => rgb <= "101001";
                when "00111000010010" => rgb <= "101001";
                when "00111000010011" => rgb <= "101001";
                when "00111000010100" => rgb <= "101001";
                when "00111000010101" => rgb <= "101000";
                when "00111000010110" => rgb <= "101001";
                when "00111000010111" => rgb <= "101001";
                when "00111000011000" => rgb <= "101001";
                when "00111000011001" => rgb <= "101001";
                when "00111000011010" => rgb <= "101000";
                when "00111000011011" => rgb <= "100100";
                when "00111000011100" => rgb <= "101000";
                when "00111000011101" => rgb <= "101000";
                when "00111000011110" => rgb <= "101000";
                when "00111000011111" => rgb <= "101000";
                when "00111000100000" => rgb <= "101000";
                when "00111000100001" => rgb <= "111001";
                when "00111000100010" => rgb <= "111001";
                when "00111000100011" => rgb <= "111001";
                when "00111000100100" => rgb <= "101001";
                when "00111000100101" => rgb <= "101000";
                when "00111000100110" => rgb <= "101000";
                when "00111000100111" => rgb <= "101001";
                when "00111000101000" => rgb <= "010000";
                when "00111000101001" => rgb <= "010000";
                when "00111000101010" => rgb <= "010000";
                when "00111000101011" => rgb <= "010000";
                when "00111010000000" => rgb <= "100001";
                when "00111010000001" => rgb <= "100001";
                when "00111010000010" => rgb <= "100001";
                when "00111010000011" => rgb <= "100101";
                when "00111010000100" => rgb <= "111010";
                when "00111010000101" => rgb <= "101001";
                when "00111010000110" => rgb <= "111001";
                when "00111010000111" => rgb <= "111001";
                when "00111010001000" => rgb <= "111001";
                when "00111010001001" => rgb <= "111001";
                when "00111010001010" => rgb <= "101001";
                when "00111010001011" => rgb <= "101001";
                when "00111010001100" => rgb <= "111001";
                when "00111010001101" => rgb <= "111001";
                when "00111010001110" => rgb <= "111001";
                when "00111010001111" => rgb <= "111001";
                when "00111010010000" => rgb <= "111001";
                when "00111010010001" => rgb <= "101001";
                when "00111010010010" => rgb <= "101001";
                when "00111010010011" => rgb <= "101001";
                when "00111010010100" => rgb <= "101000";
                when "00111010010101" => rgb <= "101000";
                when "00111010010110" => rgb <= "111001";
                when "00111010010111" => rgb <= "101001";
                when "00111010011000" => rgb <= "101001";
                when "00111010011001" => rgb <= "101001";
                when "00111010011010" => rgb <= "101000";
                when "00111010011011" => rgb <= "101000";
                when "00111010011100" => rgb <= "101000";
                when "00111010011101" => rgb <= "101000";
                when "00111010011110" => rgb <= "101000";
                when "00111010011111" => rgb <= "101000";
                when "00111010100000" => rgb <= "101000";
                when "00111010100001" => rgb <= "111001";
                when "00111010100010" => rgb <= "111001";
                when "00111010100011" => rgb <= "111001";
                when "00111010100100" => rgb <= "101001";
                when "00111010100101" => rgb <= "101000";
                when "00111010100110" => rgb <= "101000";
                when "00111010100111" => rgb <= "100100";
                when "00111010101000" => rgb <= "010000";
                when "00111010101001" => rgb <= "010000";
                when "00111010101010" => rgb <= "010000";
                when "00111010101011" => rgb <= "010000";
                when "00111100000000" => rgb <= "100001";
                when "00111100000001" => rgb <= "100001";
                when "00111100000010" => rgb <= "100001";
                when "00111100000011" => rgb <= "100101";
                when "00111100000100" => rgb <= "111010";
                when "00111100000101" => rgb <= "111001";
                when "00111100000110" => rgb <= "101001";
                when "00111100000111" => rgb <= "111001";
                when "00111100001000" => rgb <= "111001";
                when "00111100001001" => rgb <= "101001";
                when "00111100001010" => rgb <= "101001";
                when "00111100001011" => rgb <= "101001";
                when "00111100001100" => rgb <= "111001";
                when "00111100001101" => rgb <= "111001";
                when "00111100001110" => rgb <= "111001";
                when "00111100001111" => rgb <= "101001";
                when "00111100010000" => rgb <= "101001";
                when "00111100010001" => rgb <= "101001";
                when "00111100010010" => rgb <= "101001";
                when "00111100010011" => rgb <= "101001";
                when "00111100010100" => rgb <= "101000";
                when "00111100010101" => rgb <= "101000";
                when "00111100010110" => rgb <= "111001";
                when "00111100010111" => rgb <= "101001";
                when "00111100011000" => rgb <= "101001";
                when "00111100011001" => rgb <= "101001";
                when "00111100011010" => rgb <= "101000";
                when "00111100011011" => rgb <= "101000";
                when "00111100011100" => rgb <= "101000";
                when "00111100011101" => rgb <= "101000";
                when "00111100011110" => rgb <= "101000";
                when "00111100011111" => rgb <= "101000";
                when "00111100100000" => rgb <= "101000";
                when "00111100100001" => rgb <= "111001";
                when "00111100100010" => rgb <= "101001";
                when "00111100100011" => rgb <= "111001";
                when "00111100100100" => rgb <= "101001";
                when "00111100100101" => rgb <= "101000";
                when "00111100100110" => rgb <= "101000";
                when "00111100100111" => rgb <= "101000";
                when "00111100101000" => rgb <= "010000";
                when "00111100101001" => rgb <= "010000";
                when "00111100101010" => rgb <= "010000";
                when "00111100101011" => rgb <= "010000";
                when "00111110000000" => rgb <= "000000";
                when "00111110000001" => rgb <= "000000";
                when "00111110000010" => rgb <= "000000";
                when "00111110000011" => rgb <= "100101";
                when "00111110000100" => rgb <= "100101";
                when "00111110000101" => rgb <= "100101";
                when "00111110000110" => rgb <= "100101";
                when "00111110000111" => rgb <= "100101";
                when "00111110001000" => rgb <= "101001";
                when "00111110001001" => rgb <= "101001";
                when "00111110001010" => rgb <= "111001";
                when "00111110001011" => rgb <= "111001";
                when "00111110001100" => rgb <= "111001";
                when "00111110001101" => rgb <= "111001";
                when "00111110001110" => rgb <= "101001";
                when "00111110001111" => rgb <= "101001";
                when "00111110010000" => rgb <= "101001";
                when "00111110010001" => rgb <= "101001";
                when "00111110010010" => rgb <= "101001";
                when "00111110010011" => rgb <= "101001";
                when "00111110010100" => rgb <= "101000";
                when "00111110010101" => rgb <= "101000";
                when "00111110010110" => rgb <= "101001";
                when "00111110010111" => rgb <= "101001";
                when "00111110011000" => rgb <= "101001";
                when "00111110011001" => rgb <= "101000";
                when "00111110011010" => rgb <= "101000";
                when "00111110011011" => rgb <= "101000";
                when "00111110011100" => rgb <= "101000";
                when "00111110011101" => rgb <= "101001";
                when "00111110011110" => rgb <= "101001";
                when "00111110011111" => rgb <= "101001";
                when "00111110100000" => rgb <= "101001";
                when "00111110100001" => rgb <= "101001";
                when "00111110100010" => rgb <= "101001";
                when "00111110100011" => rgb <= "101001";
                when "00111110100100" => rgb <= "100101";
                when "00111110100101" => rgb <= "010100";
                when "00111110100110" => rgb <= "010000";
                when "00111110100111" => rgb <= "010000";
                when "00111110101000" => rgb <= "010000";
                when "00111110101001" => rgb <= "000000";
                when "00111110101010" => rgb <= "000000";
                when "00111110101011" => rgb <= "000000";
                when "01000000000000" => rgb <= "000000";
                when "01000000000001" => rgb <= "000000";
                when "01000000000010" => rgb <= "000000";
                when "01000000000011" => rgb <= "000000";
                when "01000000000100" => rgb <= "010001";
                when "01000000000101" => rgb <= "100001";
                when "01000000000110" => rgb <= "010001";
                when "01000000000111" => rgb <= "100101";
                when "01000000001000" => rgb <= "101001";
                when "01000000001001" => rgb <= "101001";
                when "01000000001010" => rgb <= "111001";
                when "01000000001011" => rgb <= "111001";
                when "01000000001100" => rgb <= "111001";
                when "01000000001101" => rgb <= "111001";
                when "01000000001110" => rgb <= "101001";
                when "01000000001111" => rgb <= "111001";
                when "01000000010000" => rgb <= "111001";
                when "01000000010001" => rgb <= "111001";
                when "01000000010010" => rgb <= "101001";
                when "01000000010011" => rgb <= "101001";
                when "01000000010100" => rgb <= "101000";
                when "01000000010101" => rgb <= "101000";
                when "01000000010110" => rgb <= "101000";
                when "01000000010111" => rgb <= "101000";
                when "01000000011000" => rgb <= "100100";
                when "01000000011001" => rgb <= "100100";
                when "01000000011010" => rgb <= "100100";
                when "01000000011011" => rgb <= "100100";
                when "01000000011100" => rgb <= "100100";
                when "01000000011101" => rgb <= "101001";
                when "01000000011110" => rgb <= "101001";
                when "01000000011111" => rgb <= "101001";
                when "01000000100000" => rgb <= "101001";
                when "01000000100001" => rgb <= "100100";
                when "01000000100010" => rgb <= "100100";
                when "01000000100011" => rgb <= "100100";
                when "01000000100100" => rgb <= "100100";
                when "01000000100101" => rgb <= "010000";
                when "01000000100110" => rgb <= "010000";
                when "01000000100111" => rgb <= "010000";
                when "01000000101000" => rgb <= "000000";
                when "01000000101001" => rgb <= "000000";
                when "01000000101010" => rgb <= "000000";
                when "01000000101011" => rgb <= "000000";
                when "01000010000000" => rgb <= "000000";
                when "01000010000001" => rgb <= "000000";
                when "01000010000010" => rgb <= "000000";
                when "01000010000011" => rgb <= "000000";
                when "01000010000100" => rgb <= "010001";
                when "01000010000101" => rgb <= "010001";
                when "01000010000110" => rgb <= "010001";
                when "01000010000111" => rgb <= "100101";
                when "01000010001000" => rgb <= "101001";
                when "01000010001001" => rgb <= "101001";
                when "01000010001010" => rgb <= "101001";
                when "01000010001011" => rgb <= "101001";
                when "01000010001100" => rgb <= "101001";
                when "01000010001101" => rgb <= "101001";
                when "01000010001110" => rgb <= "101001";
                when "01000010001111" => rgb <= "101001";
                when "01000010010000" => rgb <= "101001";
                when "01000010010001" => rgb <= "101001";
                when "01000010010010" => rgb <= "101001";
                when "01000010010011" => rgb <= "101001";
                when "01000010010100" => rgb <= "101000";
                when "01000010010101" => rgb <= "101000";
                when "01000010010110" => rgb <= "101000";
                when "01000010010111" => rgb <= "101000";
                when "01000010011000" => rgb <= "100100";
                when "01000010011001" => rgb <= "100100";
                when "01000010011010" => rgb <= "100100";
                when "01000010011011" => rgb <= "100100";
                when "01000010011100" => rgb <= "100100";
                when "01000010011101" => rgb <= "101001";
                when "01000010011110" => rgb <= "101001";
                when "01000010011111" => rgb <= "101001";
                when "01000010100000" => rgb <= "101001";
                when "01000010100001" => rgb <= "100100";
                when "01000010100010" => rgb <= "100100";
                when "01000010100011" => rgb <= "100100";
                when "01000010100100" => rgb <= "100100";
                when "01000010100101" => rgb <= "010000";
                when "01000010100110" => rgb <= "010000";
                when "01000010100111" => rgb <= "010000";
                when "01000010101000" => rgb <= "000000";
                when "01000010101001" => rgb <= "000000";
                when "01000010101010" => rgb <= "000000";
                when "01000010101011" => rgb <= "000000";
                when "01000100000000" => rgb <= "000000";
                when "01000100000001" => rgb <= "000000";
                when "01000100000010" => rgb <= "000000";
                when "01000100000011" => rgb <= "000000";
                when "01000100000100" => rgb <= "010001";
                when "01000100000101" => rgb <= "010001";
                when "01000100000110" => rgb <= "010001";
                when "01000100000111" => rgb <= "100101";
                when "01000100001000" => rgb <= "111001";
                when "01000100001001" => rgb <= "111001";
                when "01000100001010" => rgb <= "111001";
                when "01000100001011" => rgb <= "101001";
                when "01000100001100" => rgb <= "101001";
                when "01000100001101" => rgb <= "101001";
                when "01000100001110" => rgb <= "101001";
                when "01000100001111" => rgb <= "111001";
                when "01000100010000" => rgb <= "101001";
                when "01000100010001" => rgb <= "101001";
                when "01000100010010" => rgb <= "101001";
                when "01000100010011" => rgb <= "101001";
                when "01000100010100" => rgb <= "101001";
                when "01000100010101" => rgb <= "101000";
                when "01000100010110" => rgb <= "101000";
                when "01000100010111" => rgb <= "101000";
                when "01000100011000" => rgb <= "100100";
                when "01000100011001" => rgb <= "100100";
                when "01000100011010" => rgb <= "100100";
                when "01000100011011" => rgb <= "100100";
                when "01000100011100" => rgb <= "101000";
                when "01000100011101" => rgb <= "101001";
                when "01000100011110" => rgb <= "101001";
                when "01000100011111" => rgb <= "101001";
                when "01000100100000" => rgb <= "101001";
                when "01000100100001" => rgb <= "100100";
                when "01000100100010" => rgb <= "100100";
                when "01000100100011" => rgb <= "100100";
                when "01000100100100" => rgb <= "100100";
                when "01000100100101" => rgb <= "010000";
                when "01000100100110" => rgb <= "010000";
                when "01000100100111" => rgb <= "010000";
                when "01000100101000" => rgb <= "000000";
                when "01000100101001" => rgb <= "000000";
                when "01000100101010" => rgb <= "000000";
                when "01000100101011" => rgb <= "000000";
                when "01000110000000" => rgb <= "000000";
                when "01000110000001" => rgb <= "000000";
                when "01000110000010" => rgb <= "000000";
                when "01000110000011" => rgb <= "000000";
                when "01000110000100" => rgb <= "010001";
                when "01000110000101" => rgb <= "010001";
                when "01000110000110" => rgb <= "010001";
                when "01000110000111" => rgb <= "100101";
                when "01000110001000" => rgb <= "100101";
                when "01000110001001" => rgb <= "100101";
                when "01000110001010" => rgb <= "100101";
                when "01000110001011" => rgb <= "101001";
                when "01000110001100" => rgb <= "111001";
                when "01000110001101" => rgb <= "101001";
                when "01000110001110" => rgb <= "101001";
                when "01000110001111" => rgb <= "101001";
                when "01000110010000" => rgb <= "101001";
                when "01000110010001" => rgb <= "101001";
                when "01000110010010" => rgb <= "101001";
                when "01000110010011" => rgb <= "101001";
                when "01000110010100" => rgb <= "101001";
                when "01000110010101" => rgb <= "101000";
                when "01000110010110" => rgb <= "101001";
                when "01000110010111" => rgb <= "101001";
                when "01000110011000" => rgb <= "101001";
                when "01000110011001" => rgb <= "101001";
                when "01000110011010" => rgb <= "101001";
                when "01000110011011" => rgb <= "101001";
                when "01000110011100" => rgb <= "101001";
                when "01000110011101" => rgb <= "101000";
                when "01000110011110" => rgb <= "100100";
                when "01000110011111" => rgb <= "100100";
                when "01000110100000" => rgb <= "100100";
                when "01000110100001" => rgb <= "100100";
                when "01000110100010" => rgb <= "100100";
                when "01000110100011" => rgb <= "100100";
                when "01000110100100" => rgb <= "010000";
                when "01000110100101" => rgb <= "010000";
                when "01000110100110" => rgb <= "010000";
                when "01000110100111" => rgb <= "010000";
                when "01000110101000" => rgb <= "000000";
                when "01000110101001" => rgb <= "000000";
                when "01000110101010" => rgb <= "000000";
                when "01000110101011" => rgb <= "000000";
                when "01001000000000" => rgb <= "000000";
                when "01001000000001" => rgb <= "000000";
                when "01001000000010" => rgb <= "000000";
                when "01001000000011" => rgb <= "000000";
                when "01001000000100" => rgb <= "010001";
                when "01001000000101" => rgb <= "010001";
                when "01001000000110" => rgb <= "010001";
                when "01001000000111" => rgb <= "100101";
                when "01001000001000" => rgb <= "100101";
                when "01001000001001" => rgb <= "100101";
                when "01001000001010" => rgb <= "100101";
                when "01001000001011" => rgb <= "101001";
                when "01001000001100" => rgb <= "101001";
                when "01001000001101" => rgb <= "101001";
                when "01001000001110" => rgb <= "101001";
                when "01001000001111" => rgb <= "101001";
                when "01001000010000" => rgb <= "101001";
                when "01001000010001" => rgb <= "101001";
                when "01001000010010" => rgb <= "101001";
                when "01001000010011" => rgb <= "101001";
                when "01001000010100" => rgb <= "101001";
                when "01001000010101" => rgb <= "101000";
                when "01001000010110" => rgb <= "101001";
                when "01001000010111" => rgb <= "101001";
                when "01001000011000" => rgb <= "101001";
                when "01001000011001" => rgb <= "101001";
                when "01001000011010" => rgb <= "101001";
                when "01001000011011" => rgb <= "101001";
                when "01001000011100" => rgb <= "101001";
                when "01001000011101" => rgb <= "101000";
                when "01001000011110" => rgb <= "100100";
                when "01001000011111" => rgb <= "100100";
                when "01001000100000" => rgb <= "100100";
                when "01001000100001" => rgb <= "100100";
                when "01001000100010" => rgb <= "100100";
                when "01001000100011" => rgb <= "100100";
                when "01001000100100" => rgb <= "010000";
                when "01001000100101" => rgb <= "010000";
                when "01001000100110" => rgb <= "010000";
                when "01001000100111" => rgb <= "010000";
                when "01001000101000" => rgb <= "000000";
                when "01001000101001" => rgb <= "000000";
                when "01001000101010" => rgb <= "000000";
                when "01001000101011" => rgb <= "000000";
                when "01001010000000" => rgb <= "000000";
                when "01001010000001" => rgb <= "000000";
                when "01001010000010" => rgb <= "000000";
                when "01001010000011" => rgb <= "000000";
                when "01001010000100" => rgb <= "010001";
                when "01001010000101" => rgb <= "010001";
                when "01001010000110" => rgb <= "010001";
                when "01001010000111" => rgb <= "100101";
                when "01001010001000" => rgb <= "100101";
                when "01001010001001" => rgb <= "100101";
                when "01001010001010" => rgb <= "100101";
                when "01001010001011" => rgb <= "101001";
                when "01001010001100" => rgb <= "101001";
                when "01001010001101" => rgb <= "101001";
                when "01001010001110" => rgb <= "101001";
                when "01001010001111" => rgb <= "101001";
                when "01001010010000" => rgb <= "101001";
                when "01001010010001" => rgb <= "101001";
                when "01001010010010" => rgb <= "101001";
                when "01001010010011" => rgb <= "101001";
                when "01001010010100" => rgb <= "101001";
                when "01001010010101" => rgb <= "101000";
                when "01001010010110" => rgb <= "101001";
                when "01001010010111" => rgb <= "101001";
                when "01001010011000" => rgb <= "101001";
                when "01001010011001" => rgb <= "101001";
                when "01001010011010" => rgb <= "101001";
                when "01001010011011" => rgb <= "101001";
                when "01001010011100" => rgb <= "101001";
                when "01001010011101" => rgb <= "101000";
                when "01001010011110" => rgb <= "100100";
                when "01001010011111" => rgb <= "100100";
                when "01001010100000" => rgb <= "100100";
                when "01001010100001" => rgb <= "100100";
                when "01001010100010" => rgb <= "100100";
                when "01001010100011" => rgb <= "100100";
                when "01001010100100" => rgb <= "010000";
                when "01001010100101" => rgb <= "010000";
                when "01001010100110" => rgb <= "010000";
                when "01001010100111" => rgb <= "010000";
                when "01001010101000" => rgb <= "000000";
                when "01001010101001" => rgb <= "000000";
                when "01001010101010" => rgb <= "000000";
                when "01001010101011" => rgb <= "000000";
                when "01001100000000" => rgb <= "000000";
                when "01001100000001" => rgb <= "000000";
                when "01001100000010" => rgb <= "000000";
                when "01001100000011" => rgb <= "000000";
                when "01001100000100" => rgb <= "010001";
                when "01001100000101" => rgb <= "010001";
                when "01001100000110" => rgb <= "010001";
                when "01001100000111" => rgb <= "100101";
                when "01001100001000" => rgb <= "100101";
                when "01001100001001" => rgb <= "100101";
                when "01001100001010" => rgb <= "100101";
                when "01001100001011" => rgb <= "100101";
                when "01001100001100" => rgb <= "100101";
                when "01001100001101" => rgb <= "100101";
                when "01001100001110" => rgb <= "100101";
                when "01001100001111" => rgb <= "101001";
                when "01001100010000" => rgb <= "101001";
                when "01001100010001" => rgb <= "101001";
                when "01001100010010" => rgb <= "100101";
                when "01001100010011" => rgb <= "100101";
                when "01001100010100" => rgb <= "100101";
                when "01001100010101" => rgb <= "100100";
                when "01001100010110" => rgb <= "101001";
                when "01001100010111" => rgb <= "101001";
                when "01001100011000" => rgb <= "101001";
                when "01001100011001" => rgb <= "101001";
                when "01001100011010" => rgb <= "101000";
                when "01001100011011" => rgb <= "101000";
                when "01001100011100" => rgb <= "101000";
                when "01001100011101" => rgb <= "100100";
                when "01001100011110" => rgb <= "100100";
                when "01001100011111" => rgb <= "100100";
                when "01001100100000" => rgb <= "100100";
                when "01001100100001" => rgb <= "010100";
                when "01001100100010" => rgb <= "010100";
                when "01001100100011" => rgb <= "010100";
                when "01001100100100" => rgb <= "010000";
                when "01001100100101" => rgb <= "010000";
                when "01001100100110" => rgb <= "010000";
                when "01001100100111" => rgb <= "010000";
                when "01001100101000" => rgb <= "000000";
                when "01001100101001" => rgb <= "000000";
                when "01001100101010" => rgb <= "000000";
                when "01001100101011" => rgb <= "000000";
                when "01001110000000" => rgb <= "000000";
                when "01001110000001" => rgb <= "000000";
                when "01001110000010" => rgb <= "000000";
                when "01001110000011" => rgb <= "000000";
                when "01001110000100" => rgb <= "000000";
                when "01001110000101" => rgb <= "000000";
                when "01001110000110" => rgb <= "000000";
                when "01001110000111" => rgb <= "010001";
                when "01001110001000" => rgb <= "010001";
                when "01001110001001" => rgb <= "010001";
                when "01001110001010" => rgb <= "010001";
                when "01001110001011" => rgb <= "100101";
                when "01001110001100" => rgb <= "100101";
                when "01001110001101" => rgb <= "100101";
                when "01001110001110" => rgb <= "100101";
                when "01001110001111" => rgb <= "101001";
                when "01001110010000" => rgb <= "101001";
                when "01001110010001" => rgb <= "101001";
                when "01001110010010" => rgb <= "100101";
                when "01001110010011" => rgb <= "100101";
                when "01001110010100" => rgb <= "100100";
                when "01001110010101" => rgb <= "100100";
                when "01001110010110" => rgb <= "100100";
                when "01001110010111" => rgb <= "100100";
                when "01001110011000" => rgb <= "100100";
                when "01001110011001" => rgb <= "100100";
                when "01001110011010" => rgb <= "100100";
                when "01001110011011" => rgb <= "100100";
                when "01001110011100" => rgb <= "100100";
                when "01001110011101" => rgb <= "100100";
                when "01001110011110" => rgb <= "100100";
                when "01001110011111" => rgb <= "100100";
                when "01001110100000" => rgb <= "100100";
                when "01001110100001" => rgb <= "010000";
                when "01001110100010" => rgb <= "010000";
                when "01001110100011" => rgb <= "010000";
                when "01001110100100" => rgb <= "000000";
                when "01001110100101" => rgb <= "000000";
                when "01001110100110" => rgb <= "000000";
                when "01001110100111" => rgb <= "000000";
                when "01001110101000" => rgb <= "000000";
                when "01001110101001" => rgb <= "000000";
                when "01001110101010" => rgb <= "000000";
                when "01001110101011" => rgb <= "000000";
                when "01010000000000" => rgb <= "000000";
                when "01010000000001" => rgb <= "000000";
                when "01010000000010" => rgb <= "000000";
                when "01010000000011" => rgb <= "000000";
                when "01010000000100" => rgb <= "000000";
                when "01010000000101" => rgb <= "000000";
                when "01010000000110" => rgb <= "000000";
                when "01010000000111" => rgb <= "010001";
                when "01010000001000" => rgb <= "010001";
                when "01010000001001" => rgb <= "010001";
                when "01010000001010" => rgb <= "010001";
                when "01010000001011" => rgb <= "100101";
                when "01010000001100" => rgb <= "100101";
                when "01010000001101" => rgb <= "100101";
                when "01010000001110" => rgb <= "100101";
                when "01010000001111" => rgb <= "101001";
                when "01010000010000" => rgb <= "101001";
                when "01010000010001" => rgb <= "101001";
                when "01010000010010" => rgb <= "100101";
                when "01010000010011" => rgb <= "100101";
                when "01010000010100" => rgb <= "100100";
                when "01010000010101" => rgb <= "100100";
                when "01010000010110" => rgb <= "100100";
                when "01010000010111" => rgb <= "100100";
                when "01010000011000" => rgb <= "100100";
                when "01010000011001" => rgb <= "100100";
                when "01010000011010" => rgb <= "100100";
                when "01010000011011" => rgb <= "100100";
                when "01010000011100" => rgb <= "100100";
                when "01010000011101" => rgb <= "100100";
                when "01010000011110" => rgb <= "100100";
                when "01010000011111" => rgb <= "100100";
                when "01010000100000" => rgb <= "100100";
                when "01010000100001" => rgb <= "010000";
                when "01010000100010" => rgb <= "010000";
                when "01010000100011" => rgb <= "010000";
                when "01010000100100" => rgb <= "000000";
                when "01010000100101" => rgb <= "000000";
                when "01010000100110" => rgb <= "000000";
                when "01010000100111" => rgb <= "000000";
                when "01010000101000" => rgb <= "000000";
                when "01010000101001" => rgb <= "000000";
                when "01010000101010" => rgb <= "000000";
                when "01010000101011" => rgb <= "000000";
                when "01010010000000" => rgb <= "000000";
                when "01010010000001" => rgb <= "000000";
                when "01010010000010" => rgb <= "000000";
                when "01010010000011" => rgb <= "000000";
                when "01010010000100" => rgb <= "000000";
                when "01010010000101" => rgb <= "000000";
                when "01010010000110" => rgb <= "000000";
                when "01010010000111" => rgb <= "010001";
                when "01010010001000" => rgb <= "010001";
                when "01010010001001" => rgb <= "010001";
                when "01010010001010" => rgb <= "010001";
                when "01010010001011" => rgb <= "100101";
                when "01010010001100" => rgb <= "100101";
                when "01010010001101" => rgb <= "100101";
                when "01010010001110" => rgb <= "100101";
                when "01010010001111" => rgb <= "101001";
                when "01010010010000" => rgb <= "101001";
                when "01010010010001" => rgb <= "101001";
                when "01010010010010" => rgb <= "100101";
                when "01010010010011" => rgb <= "100101";
                when "01010010010100" => rgb <= "100100";
                when "01010010010101" => rgb <= "100100";
                when "01010010010110" => rgb <= "100100";
                when "01010010010111" => rgb <= "100100";
                when "01010010011000" => rgb <= "100100";
                when "01010010011001" => rgb <= "100100";
                when "01010010011010" => rgb <= "100100";
                when "01010010011011" => rgb <= "100100";
                when "01010010011100" => rgb <= "100100";
                when "01010010011101" => rgb <= "100100";
                when "01010010011110" => rgb <= "100100";
                when "01010010011111" => rgb <= "100100";
                when "01010010100000" => rgb <= "100100";
                when "01010010100001" => rgb <= "010000";
                when "01010010100010" => rgb <= "010000";
                when "01010010100011" => rgb <= "010000";
                when "01010010100100" => rgb <= "000000";
                when "01010010100101" => rgb <= "000000";
                when "01010010100110" => rgb <= "000000";
                when "01010010100111" => rgb <= "000000";
                when "01010010101000" => rgb <= "000000";
                when "01010010101001" => rgb <= "000000";
                when "01010010101010" => rgb <= "000000";
                when "01010010101011" => rgb <= "000000";
                when "01010100000000" => rgb <= "000000";
                when "01010100000001" => rgb <= "000000";
                when "01010100000010" => rgb <= "000000";
                when "01010100000011" => rgb <= "000000";
                when "01010100000100" => rgb <= "000000";
                when "01010100000101" => rgb <= "000000";
                when "01010100000110" => rgb <= "000000";
                when "01010100000111" => rgb <= "000000";
                when "01010100001000" => rgb <= "000000";
                when "01010100001001" => rgb <= "000000";
                when "01010100001010" => rgb <= "000000";
                when "01010100001011" => rgb <= "010001";
                when "01010100001100" => rgb <= "010001";
                when "01010100001101" => rgb <= "010001";
                when "01010100001110" => rgb <= "010001";
                when "01010100001111" => rgb <= "100101";
                when "01010100010000" => rgb <= "100100";
                when "01010100010001" => rgb <= "100100";
                when "01010100010010" => rgb <= "010000";
                when "01010100010011" => rgb <= "010000";
                when "01010100010100" => rgb <= "010000";
                when "01010100010101" => rgb <= "010000";
                when "01010100010110" => rgb <= "010000";
                when "01010100010111" => rgb <= "010000";
                when "01010100011000" => rgb <= "010000";
                when "01010100011001" => rgb <= "010000";
                when "01010100011010" => rgb <= "010000";
                when "01010100011011" => rgb <= "010000";
                when "01010100011100" => rgb <= "010000";
                when "01010100011101" => rgb <= "010000";
                when "01010100011110" => rgb <= "010000";
                when "01010100011111" => rgb <= "010000";
                when "01010100100000" => rgb <= "010000";
                when "01010100100001" => rgb <= "000000";
                when "01010100100010" => rgb <= "000000";
                when "01010100100011" => rgb <= "000000";
                when "01010100100100" => rgb <= "000000";
                when "01010100100101" => rgb <= "000000";
                when "01010100100110" => rgb <= "000000";
                when "01010100100111" => rgb <= "000000";
                when "01010100101000" => rgb <= "000000";
                when "01010100101001" => rgb <= "000000";
                when "01010100101010" => rgb <= "000000";
                when "01010100101011" => rgb <= "000000";
                when "01010110000000" => rgb <= "000000";
                when "01010110000001" => rgb <= "000000";
                when "01010110000010" => rgb <= "000000";
                when "01010110000011" => rgb <= "000000";
                when "01010110000100" => rgb <= "000000";
                when "01010110000101" => rgb <= "000000";
                when "01010110000110" => rgb <= "000000";
                when "01010110000111" => rgb <= "000000";
                when "01010110001000" => rgb <= "000000";
                when "01010110001001" => rgb <= "000000";
                when "01010110001010" => rgb <= "000000";
                when "01010110001011" => rgb <= "010001";
                when "01010110001100" => rgb <= "010001";
                when "01010110001101" => rgb <= "010001";
                when "01010110001110" => rgb <= "010000";
                when "01010110001111" => rgb <= "010000";
                when "01010110010000" => rgb <= "010000";
                when "01010110010001" => rgb <= "010000";
                when "01010110010010" => rgb <= "010000";
                when "01010110010011" => rgb <= "010000";
                when "01010110010100" => rgb <= "010000";
                when "01010110010101" => rgb <= "010000";
                when "01010110010110" => rgb <= "010000";
                when "01010110010111" => rgb <= "010000";
                when "01010110011000" => rgb <= "010000";
                when "01010110011001" => rgb <= "010000";
                when "01010110011010" => rgb <= "010000";
                when "01010110011011" => rgb <= "010000";
                when "01010110011100" => rgb <= "010000";
                when "01010110011101" => rgb <= "010000";
                when "01010110011110" => rgb <= "010000";
                when "01010110011111" => rgb <= "010000";
                when "01010110100000" => rgb <= "010000";
                when "01010110100001" => rgb <= "000000";
                when "01010110100010" => rgb <= "000000";
                when "01010110100011" => rgb <= "000000";
                when "01010110100100" => rgb <= "000000";
                when "01010110100101" => rgb <= "000000";
                when "01010110100110" => rgb <= "000000";
                when "01010110100111" => rgb <= "000000";
                when "01010110101000" => rgb <= "000000";
                when "01010110101001" => rgb <= "000000";
                when "01010110101010" => rgb <= "000000";
                when "01010110101011" => rgb <= "000000";
                when others => rgb <= "111111";
               
                end case;
            end if;
            end process;
        end;
                
