library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity one_segments is
    port (
        row : in unsigned (9 downto 0);
        col : in unsigned (9 downto 0);
        clk : in std_logic;
        rgb : out std_logic_vector(5 downto 0)
    );
end one_segments;

architecture synth of one_segments is
    signal addr : std_logic_vector(13 downto 0);

    begin
        addr <= std_logic_vector(row(7 downto 0)) & std_logic_vector(col(7 downto 0));
        process(clk) is begin
            if rising_edge(clk) then 
                case addr is 
                when "00000000000000" => rgb <= "000000";
                when "00000000000001" => rgb <= "000000";
                when "00000000000010" => rgb <= "000000";
                when "00000000000011" => rgb <= "000000";
                when "00000000000100" => rgb <= "000000";
                when "00000000000101" => rgb <= "000000";
                when "00000000000110" => rgb <= "000000";
                when "00000000000111" => rgb <= "000000";
                when "00000000001000" => rgb <= "000000";
                when "00000000001001" => rgb <= "000000";
                when "00000000001010" => rgb <= "000000";
                when "00000000001011" => rgb <= "000000";
                when "00000000001100" => rgb <= "000000";
                when "00000000001101" => rgb <= "000000";
                when "00000000001110" => rgb <= "000000";
                when "00000000001111" => rgb <= "000000";
                when "00000000010000" => rgb <= "000000";
                when "00000000010001" => rgb <= "000000";
                when "00000000010010" => rgb <= "000000";
                when "00000000010011" => rgb <= "000000";
                when "00000000010100" => rgb <= "000000";
                when "00000000010101" => rgb <= "000000";
                when "00000000010110" => rgb <= "000000";
                when "00000000010111" => rgb <= "000000";
                when "00000000011000" => rgb <= "000000";
                when "00000000011001" => rgb <= "000000";
                when "00000000011010" => rgb <= "000000";
                when "00000000011011" => rgb <= "000000";
                when "00000000011100" => rgb <= "000000";
                when "00000000011101" => rgb <= "000000";
                when "00000000011110" => rgb <= "000000";
                when "00000000011111" => rgb <= "000011";
                when "00000000100000" => rgb <= "000011";
                when "00000000100001" => rgb <= "000011";
                when "00000000100010" => rgb <= "000011";
                when "00000010000000" => rgb <= "000000";
                when "00000010000001" => rgb <= "000000";
                when "00000010000010" => rgb <= "000000";
                when "00000010000011" => rgb <= "000000";
                when "00000010000100" => rgb <= "000000";
                when "00000010000101" => rgb <= "000000";
                when "00000010000110" => rgb <= "000000";
                when "00000010000111" => rgb <= "000000";
                when "00000010001000" => rgb <= "000000";
                when "00000010001001" => rgb <= "000000";
                when "00000010001010" => rgb <= "000000";
                when "00000010001011" => rgb <= "000000";
                when "00000010001100" => rgb <= "000000";
                when "00000010001101" => rgb <= "000000";
                when "00000010001110" => rgb <= "000000";
                when "00000010001111" => rgb <= "000000";
                when "00000010010000" => rgb <= "000000";
                when "00000010010001" => rgb <= "000000";
                when "00000010010010" => rgb <= "000000";
                when "00000010010011" => rgb <= "000000";
                when "00000010010100" => rgb <= "000000";
                when "00000010010101" => rgb <= "000000";
                when "00000010010110" => rgb <= "000000";
                when "00000010010111" => rgb <= "000000";
                when "00000010011000" => rgb <= "000000";
                when "00000010011001" => rgb <= "000000";
                when "00000010011010" => rgb <= "000000";
                when "00000010011011" => rgb <= "000000";
                when "00000010011100" => rgb <= "000000";
                when "00000010011101" => rgb <= "000000";
                when "00000010011110" => rgb <= "000000";
                when "00000010011111" => rgb <= "000011";
                when "00000010100000" => rgb <= "000011";
                when "00000010100001" => rgb <= "000011";
                when "00000010100010" => rgb <= "000011";
                when "00000100000000" => rgb <= "000000";
                when "00000100000001" => rgb <= "000000";
                when "00000100000010" => rgb <= "000000";
                when "00000100000011" => rgb <= "000000";
                when "00000100000100" => rgb <= "000000";
                when "00000100000101" => rgb <= "000000";
                when "00000100000110" => rgb <= "000000";
                when "00000100000111" => rgb <= "000000";
                when "00000100001000" => rgb <= "000000";
                when "00000100001001" => rgb <= "000000";
                when "00000100001010" => rgb <= "000000";
                when "00000100001011" => rgb <= "000000";
                when "00000100001100" => rgb <= "000000";
                when "00000100001101" => rgb <= "000000";
                when "00000100001110" => rgb <= "000000";
                when "00000100001111" => rgb <= "000000";
                when "00000100010000" => rgb <= "000000";
                when "00000100010001" => rgb <= "000000";
                when "00000100010010" => rgb <= "000000";
                when "00000100010011" => rgb <= "000000";
                when "00000100010100" => rgb <= "000000";
                when "00000100010101" => rgb <= "000000";
                when "00000100010110" => rgb <= "000000";
                when "00000100010111" => rgb <= "000000";
                when "00000100011000" => rgb <= "000000";
                when "00000100011001" => rgb <= "000000";
                when "00000100011010" => rgb <= "000000";
                when "00000100011011" => rgb <= "000000";
                when "00000100011100" => rgb <= "000000";
                when "00000100011101" => rgb <= "000000";
                when "00000100011110" => rgb <= "000000";
                when "00000100011111" => rgb <= "000011";
                when "00000100100000" => rgb <= "000011";
                when "00000100100001" => rgb <= "000011";
                when "00000100100010" => rgb <= "000011";
                when "00000110000000" => rgb <= "000000";
                when "00000110000001" => rgb <= "000000";
                when "00000110000010" => rgb <= "000000";
                when "00000110000011" => rgb <= "000000";
                when "00000110000100" => rgb <= "000000";
                when "00000110000101" => rgb <= "000000";
                when "00000110000110" => rgb <= "000000";
                when "00000110000111" => rgb <= "000000";
                when "00000110001000" => rgb <= "000000";
                when "00000110001001" => rgb <= "000000";
                when "00000110001010" => rgb <= "000000";
                when "00000110001011" => rgb <= "000000";
                when "00000110001100" => rgb <= "000000";
                when "00000110001101" => rgb <= "000000";
                when "00000110001110" => rgb <= "000000";
                when "00000110001111" => rgb <= "000000";
                when "00000110010000" => rgb <= "000000";
                when "00000110010001" => rgb <= "000000";
                when "00000110010010" => rgb <= "000000";
                when "00000110010011" => rgb <= "000000";
                when "00000110010100" => rgb <= "000000";
                when "00000110010101" => rgb <= "000000";
                when "00000110010110" => rgb <= "000000";
                when "00000110010111" => rgb <= "000000";
                when "00000110011000" => rgb <= "000000";
                when "00000110011001" => rgb <= "000000";
                when "00000110011010" => rgb <= "000000";
                when "00000110011011" => rgb <= "000000";
                when "00000110011100" => rgb <= "000000";
                when "00000110011101" => rgb <= "000000";
                when "00000110011110" => rgb <= "000000";
                when "00000110011111" => rgb <= "000011";
                when "00000110100000" => rgb <= "000011";
                when "00000110100001" => rgb <= "000011";
                when "00000110100010" => rgb <= "000011";
                when "00001000000000" => rgb <= "000000";
                when "00001000000001" => rgb <= "000000";
                when "00001000000010" => rgb <= "000000";
                when "00001000000011" => rgb <= "000000";
                when "00001000000100" => rgb <= "000000";
                when "00001000000101" => rgb <= "000000";
                when "00001000000110" => rgb <= "000000";
                when "00001000000111" => rgb <= "000000";
                when "00001000001000" => rgb <= "000000";
                when "00001000001001" => rgb <= "000000";
                when "00001000001010" => rgb <= "000000";
                when "00001000001011" => rgb <= "000000";
                when "00001000001100" => rgb <= "000000";
                when "00001000001101" => rgb <= "000000";
                when "00001000001110" => rgb <= "000000";
                when "00001000001111" => rgb <= "000000";
                when "00001000010000" => rgb <= "000000";
                when "00001000010001" => rgb <= "000000";
                when "00001000010010" => rgb <= "000000";
                when "00001000010011" => rgb <= "000000";
                when "00001000010100" => rgb <= "000000";
                when "00001000010101" => rgb <= "000000";
                when "00001000010110" => rgb <= "000000";
                when "00001000010111" => rgb <= "000000";
                when "00001000011000" => rgb <= "000000";
                when "00001000011001" => rgb <= "000000";
                when "00001000011010" => rgb <= "000000";
                when "00001000011011" => rgb <= "000000";
                when "00001000011100" => rgb <= "000000";
                when "00001000011101" => rgb <= "000000";
                when "00001000011110" => rgb <= "000000";
                when "00001000011111" => rgb <= "000011";
                when "00001000100000" => rgb <= "000011";
                when "00001000100001" => rgb <= "000011";
                when "00001000100010" => rgb <= "000011";
                when "00001010000000" => rgb <= "000000";
                when "00001010000001" => rgb <= "000000";
                when "00001010000010" => rgb <= "000000";
                when "00001010000011" => rgb <= "000000";
                when "00001010000100" => rgb <= "000000";
                when "00001010000101" => rgb <= "000000";
                when "00001010000110" => rgb <= "000000";
                when "00001010000111" => rgb <= "000000";
                when "00001010001000" => rgb <= "000000";
                when "00001010001001" => rgb <= "000000";
                when "00001010001010" => rgb <= "000000";
                when "00001010001011" => rgb <= "000000";
                when "00001010001100" => rgb <= "000000";
                when "00001010001101" => rgb <= "000000";
                when "00001010001110" => rgb <= "000000";
                when "00001010001111" => rgb <= "000000";
                when "00001010010000" => rgb <= "000000";
                when "00001010010001" => rgb <= "000000";
                when "00001010010010" => rgb <= "000000";
                when "00001010010011" => rgb <= "000000";
                when "00001010010100" => rgb <= "000000";
                when "00001010010101" => rgb <= "000000";
                when "00001010010110" => rgb <= "000000";
                when "00001010010111" => rgb <= "000000";
                when "00001010011000" => rgb <= "000000";
                when "00001010011001" => rgb <= "000000";
                when "00001010011010" => rgb <= "000000";
                when "00001010011011" => rgb <= "000000";
                when "00001010011100" => rgb <= "000000";
                when "00001010011101" => rgb <= "000000";
                when "00001010011110" => rgb <= "000000";
                when "00001010011111" => rgb <= "000011";
                when "00001010100000" => rgb <= "000011";
                when "00001010100001" => rgb <= "000011";
                when "00001010100010" => rgb <= "000011";
                when "00001100000000" => rgb <= "000000";
                when "00001100000001" => rgb <= "000000";
                when "00001100000010" => rgb <= "000000";
                when "00001100000011" => rgb <= "000000";
                when "00001100000100" => rgb <= "000000";
                when "00001100000101" => rgb <= "000000";
                when "00001100000110" => rgb <= "000000";
                when "00001100000111" => rgb <= "000000";
                when "00001100001000" => rgb <= "000000";
                when "00001100001001" => rgb <= "000000";
                when "00001100001010" => rgb <= "000000";
                when "00001100001011" => rgb <= "000000";
                when "00001100001100" => rgb <= "000000";
                when "00001100001101" => rgb <= "000000";
                when "00001100001110" => rgb <= "000000";
                when "00001100001111" => rgb <= "000000";
                when "00001100010000" => rgb <= "000000";
                when "00001100010001" => rgb <= "000000";
                when "00001100010010" => rgb <= "000000";
                when "00001100010011" => rgb <= "000000";
                when "00001100010100" => rgb <= "000000";
                when "00001100010101" => rgb <= "000000";
                when "00001100010110" => rgb <= "000000";
                when "00001100010111" => rgb <= "000000";
                when "00001100011000" => rgb <= "000000";
                when "00001100011001" => rgb <= "000000";
                when "00001100011010" => rgb <= "000000";
                when "00001100011011" => rgb <= "000000";
                when "00001100011100" => rgb <= "000000";
                when "00001100011101" => rgb <= "000000";
                when "00001100011110" => rgb <= "000000";
                when "00001100011111" => rgb <= "000011";
                when "00001100100000" => rgb <= "000011";
                when "00001100100001" => rgb <= "000011";
                when "00001100100010" => rgb <= "000011";
                when "00001110000000" => rgb <= "000000";
                when "00001110000001" => rgb <= "000000";
                when "00001110000010" => rgb <= "000000";
                when "00001110000011" => rgb <= "000000";
                when "00001110000100" => rgb <= "000000";
                when "00001110000101" => rgb <= "000000";
                when "00001110000110" => rgb <= "000000";
                when "00001110000111" => rgb <= "000000";
                when "00001110001000" => rgb <= "000000";
                when "00001110001001" => rgb <= "000000";
                when "00001110001010" => rgb <= "000000";
                when "00001110001011" => rgb <= "000000";
                when "00001110001100" => rgb <= "000000";
                when "00001110001101" => rgb <= "000000";
                when "00001110001110" => rgb <= "000000";
                when "00001110001111" => rgb <= "000000";
                when "00001110010000" => rgb <= "000000";
                when "00001110010001" => rgb <= "000000";
                when "00001110010010" => rgb <= "000000";
                when "00001110010011" => rgb <= "000000";
                when "00001110010100" => rgb <= "000000";
                when "00001110010101" => rgb <= "000000";
                when "00001110010110" => rgb <= "000000";
                when "00001110010111" => rgb <= "000000";
                when "00001110011000" => rgb <= "000000";
                when "00001110011001" => rgb <= "000000";
                when "00001110011010" => rgb <= "000000";
                when "00001110011011" => rgb <= "000000";
                when "00001110011100" => rgb <= "000000";
                when "00001110011101" => rgb <= "000000";
                when "00001110011110" => rgb <= "000000";
                when "00001110011111" => rgb <= "000011";
                when "00001110100000" => rgb <= "000011";
                when "00001110100001" => rgb <= "000011";
                when "00001110100010" => rgb <= "000011";
                when "00010000000000" => rgb <= "000000";
                when "00010000000001" => rgb <= "000000";
                when "00010000000010" => rgb <= "000000";
                when "00010000000011" => rgb <= "000000";
                when "00010000000100" => rgb <= "000000";
                when "00010000000101" => rgb <= "000000";
                when "00010000000110" => rgb <= "000000";
                when "00010000000111" => rgb <= "000000";
                when "00010000001000" => rgb <= "000000";
                when "00010000001001" => rgb <= "000000";
                when "00010000001010" => rgb <= "000000";
                when "00010000001011" => rgb <= "000000";
                when "00010000001100" => rgb <= "000000";
                when "00010000001101" => rgb <= "000000";
                when "00010000001110" => rgb <= "000000";
                when "00010000001111" => rgb <= "000000";
                when "00010000010000" => rgb <= "000000";
                when "00010000010001" => rgb <= "000000";
                when "00010000010010" => rgb <= "000000";
                when "00010000010011" => rgb <= "000000";
                when "00010000010100" => rgb <= "000000";
                when "00010000010101" => rgb <= "000000";
                when "00010000010110" => rgb <= "000000";
                when "00010000010111" => rgb <= "000000";
                when "00010000011000" => rgb <= "000000";
                when "00010000011001" => rgb <= "000000";
                when "00010000011010" => rgb <= "000000";
                when "00010000011011" => rgb <= "000000";
                when "00010000011100" => rgb <= "000000";
                when "00010000011101" => rgb <= "000000";
                when "00010000011110" => rgb <= "000000";
                when "00010000011111" => rgb <= "000011";
                when "00010000100000" => rgb <= "000011";
                when "00010000100001" => rgb <= "000011";
                when "00010000100010" => rgb <= "000011";
                when "00010010000000" => rgb <= "000000";
                when "00010010000001" => rgb <= "000000";
                when "00010010000010" => rgb <= "000000";
                when "00010010000011" => rgb <= "000000";
                when "00010010000100" => rgb <= "000000";
                when "00010010000101" => rgb <= "000000";
                when "00010010000110" => rgb <= "000000";
                when "00010010000111" => rgb <= "000000";
                when "00010010001000" => rgb <= "000000";
                when "00010010001001" => rgb <= "000000";
                when "00010010001010" => rgb <= "000000";
                when "00010010001011" => rgb <= "000000";
                when "00010010001100" => rgb <= "000000";
                when "00010010001101" => rgb <= "000000";
                when "00010010001110" => rgb <= "000000";
                when "00010010001111" => rgb <= "000000";
                when "00010010010000" => rgb <= "000000";
                when "00010010010001" => rgb <= "000000";
                when "00010010010010" => rgb <= "000000";
                when "00010010010011" => rgb <= "000000";
                when "00010010010100" => rgb <= "000000";
                when "00010010010101" => rgb <= "000000";
                when "00010010010110" => rgb <= "000000";
                when "00010010010111" => rgb <= "000000";
                when "00010010011000" => rgb <= "000000";
                when "00010010011001" => rgb <= "000000";
                when "00010010011010" => rgb <= "000000";
                when "00010010011011" => rgb <= "000000";
                when "00010010011100" => rgb <= "000000";
                when "00010010011101" => rgb <= "000000";
                when "00010010011110" => rgb <= "000000";
                when "00010010011111" => rgb <= "000011";
                when "00010010100000" => rgb <= "000011";
                when "00010010100001" => rgb <= "000011";
                when "00010010100010" => rgb <= "000011";
                when "00010100000000" => rgb <= "000000";
                when "00010100000001" => rgb <= "000000";
                when "00010100000010" => rgb <= "000000";
                when "00010100000011" => rgb <= "000000";
                when "00010100000100" => rgb <= "000000";
                when "00010100000101" => rgb <= "000000";
                when "00010100000110" => rgb <= "000000";
                when "00010100000111" => rgb <= "000000";
                when "00010100001000" => rgb <= "000000";
                when "00010100001001" => rgb <= "000000";
                when "00010100001010" => rgb <= "000000";
                when "00010100001011" => rgb <= "000000";
                when "00010100001100" => rgb <= "000000";
                when "00010100001101" => rgb <= "000000";
                when "00010100001110" => rgb <= "000000";
                when "00010100001111" => rgb <= "000000";
                when "00010100010000" => rgb <= "000000";
                when "00010100010001" => rgb <= "000000";
                when "00010100010010" => rgb <= "000000";
                when "00010100010011" => rgb <= "000000";
                when "00010100010100" => rgb <= "000000";
                when "00010100010101" => rgb <= "000000";
                when "00010100010110" => rgb <= "000000";
                when "00010100010111" => rgb <= "000000";
                when "00010100011000" => rgb <= "000000";
                when "00010100011001" => rgb <= "000000";
                when "00010100011010" => rgb <= "000000";
                when "00010100011011" => rgb <= "000000";
                when "00010100011100" => rgb <= "000000";
                when "00010100011101" => rgb <= "000000";
                when "00010100011110" => rgb <= "000000";
                when "00010100011111" => rgb <= "000011";
                when "00010100100000" => rgb <= "000011";
                when "00010100100001" => rgb <= "000011";
                when "00010100100010" => rgb <= "000011";
                when "00010110000000" => rgb <= "000000";
                when "00010110000001" => rgb <= "000000";
                when "00010110000010" => rgb <= "000000";
                when "00010110000011" => rgb <= "000000";
                when "00010110000100" => rgb <= "000000";
                when "00010110000101" => rgb <= "000000";
                when "00010110000110" => rgb <= "000000";
                when "00010110000111" => rgb <= "000000";
                when "00010110001000" => rgb <= "000000";
                when "00010110001001" => rgb <= "000000";
                when "00010110001010" => rgb <= "000000";
                when "00010110001011" => rgb <= "000000";
                when "00010110001100" => rgb <= "000000";
                when "00010110001101" => rgb <= "000000";
                when "00010110001110" => rgb <= "000000";
                when "00010110001111" => rgb <= "000000";
                when "00010110010000" => rgb <= "000000";
                when "00010110010001" => rgb <= "000000";
                when "00010110010010" => rgb <= "000000";
                when "00010110010011" => rgb <= "000000";
                when "00010110010100" => rgb <= "000000";
                when "00010110010101" => rgb <= "000000";
                when "00010110010110" => rgb <= "000000";
                when "00010110010111" => rgb <= "000000";
                when "00010110011000" => rgb <= "000000";
                when "00010110011001" => rgb <= "000000";
                when "00010110011010" => rgb <= "000000";
                when "00010110011011" => rgb <= "000000";
                when "00010110011100" => rgb <= "000000";
                when "00010110011101" => rgb <= "000000";
                when "00010110011110" => rgb <= "000000";
                when "00010110011111" => rgb <= "000011";
                when "00010110100000" => rgb <= "000011";
                when "00010110100001" => rgb <= "000011";
                when "00010110100010" => rgb <= "000011";
                when "00011000000000" => rgb <= "000000";
                when "00011000000001" => rgb <= "000000";
                when "00011000000010" => rgb <= "000000";
                when "00011000000011" => rgb <= "000000";
                when "00011000000100" => rgb <= "000000";
                when "00011000000101" => rgb <= "000000";
                when "00011000000110" => rgb <= "000000";
                when "00011000000111" => rgb <= "000000";
                when "00011000001000" => rgb <= "000000";
                when "00011000001001" => rgb <= "000000";
                when "00011000001010" => rgb <= "000000";
                when "00011000001011" => rgb <= "000000";
                when "00011000001100" => rgb <= "000000";
                when "00011000001101" => rgb <= "000000";
                when "00011000001110" => rgb <= "000000";
                when "00011000001111" => rgb <= "000000";
                when "00011000010000" => rgb <= "000000";
                when "00011000010001" => rgb <= "000000";
                when "00011000010010" => rgb <= "000000";
                when "00011000010011" => rgb <= "000000";
                when "00011000010100" => rgb <= "000000";
                when "00011000010101" => rgb <= "000000";
                when "00011000010110" => rgb <= "000000";
                when "00011000010111" => rgb <= "000000";
                when "00011000011000" => rgb <= "000000";
                when "00011000011001" => rgb <= "000000";
                when "00011000011010" => rgb <= "000000";
                when "00011000011011" => rgb <= "000000";
                when "00011000011100" => rgb <= "000000";
                when "00011000011101" => rgb <= "000000";
                when "00011000011110" => rgb <= "000000";
                when "00011000011111" => rgb <= "000011";
                when "00011000100000" => rgb <= "000011";
                when "00011000100001" => rgb <= "000011";
                when "00011000100010" => rgb <= "000011";
                when "00011010000000" => rgb <= "000000";
                when "00011010000001" => rgb <= "000000";
                when "00011010000010" => rgb <= "000000";
                when "00011010000011" => rgb <= "000000";
                when "00011010000100" => rgb <= "000000";
                when "00011010000101" => rgb <= "000000";
                when "00011010000110" => rgb <= "000000";
                when "00011010000111" => rgb <= "000000";
                when "00011010001000" => rgb <= "000000";
                when "00011010001001" => rgb <= "000000";
                when "00011010001010" => rgb <= "000000";
                when "00011010001011" => rgb <= "000000";
                when "00011010001100" => rgb <= "000000";
                when "00011010001101" => rgb <= "000000";
                when "00011010001110" => rgb <= "000000";
                when "00011010001111" => rgb <= "000000";
                when "00011010010000" => rgb <= "000000";
                when "00011010010001" => rgb <= "000000";
                when "00011010010010" => rgb <= "000000";
                when "00011010010011" => rgb <= "000000";
                when "00011010010100" => rgb <= "000000";
                when "00011010010101" => rgb <= "000000";
                when "00011010010110" => rgb <= "000000";
                when "00011010010111" => rgb <= "000000";
                when "00011010011000" => rgb <= "000000";
                when "00011010011001" => rgb <= "000000";
                when "00011010011010" => rgb <= "000000";
                when "00011010011011" => rgb <= "000000";
                when "00011010011100" => rgb <= "000000";
                when "00011010011101" => rgb <= "000000";
                when "00011010011110" => rgb <= "000000";
                when "00011010011111" => rgb <= "000011";
                when "00011010100000" => rgb <= "000011";
                when "00011010100001" => rgb <= "000011";
                when "00011010100010" => rgb <= "000011";
                when "00011100000000" => rgb <= "000000";
                when "00011100000001" => rgb <= "000000";
                when "00011100000010" => rgb <= "000000";
                when "00011100000011" => rgb <= "000000";
                when "00011100000100" => rgb <= "000000";
                when "00011100000101" => rgb <= "000000";
                when "00011100000110" => rgb <= "000000";
                when "00011100000111" => rgb <= "000000";
                when "00011100001000" => rgb <= "000000";
                when "00011100001001" => rgb <= "000000";
                when "00011100001010" => rgb <= "000000";
                when "00011100001011" => rgb <= "000000";
                when "00011100001100" => rgb <= "000000";
                when "00011100001101" => rgb <= "000000";
                when "00011100001110" => rgb <= "000000";
                when "00011100001111" => rgb <= "000000";
                when "00011100010000" => rgb <= "000000";
                when "00011100010001" => rgb <= "000000";
                when "00011100010010" => rgb <= "000000";
                when "00011100010011" => rgb <= "000000";
                when "00011100010100" => rgb <= "000000";
                when "00011100010101" => rgb <= "000000";
                when "00011100010110" => rgb <= "000000";
                when "00011100010111" => rgb <= "000000";
                when "00011100011000" => rgb <= "000000";
                when "00011100011001" => rgb <= "000000";
                when "00011100011010" => rgb <= "000000";
                when "00011100011011" => rgb <= "000000";
                when "00011100011100" => rgb <= "000000";
                when "00011100011101" => rgb <= "000000";
                when "00011100011110" => rgb <= "000000";
                when "00011100011111" => rgb <= "000011";
                when "00011100100000" => rgb <= "000011";
                when "00011100100001" => rgb <= "000011";
                when "00011100100010" => rgb <= "000011";
                when "00011110000000" => rgb <= "000000";
                when "00011110000001" => rgb <= "000000";
                when "00011110000010" => rgb <= "000000";
                when "00011110000011" => rgb <= "000000";
                when "00011110000100" => rgb <= "000000";
                when "00011110000101" => rgb <= "000000";
                when "00011110000110" => rgb <= "000000";
                when "00011110000111" => rgb <= "000000";
                when "00011110001000" => rgb <= "000000";
                when "00011110001001" => rgb <= "000000";
                when "00011110001010" => rgb <= "000000";
                when "00011110001011" => rgb <= "000000";
                when "00011110001100" => rgb <= "000000";
                when "00011110001101" => rgb <= "000000";
                when "00011110001110" => rgb <= "000000";
                when "00011110001111" => rgb <= "000000";
                when "00011110010000" => rgb <= "000000";
                when "00011110010001" => rgb <= "000000";
                when "00011110010010" => rgb <= "000000";
                when "00011110010011" => rgb <= "000000";
                when "00011110010100" => rgb <= "000000";
                when "00011110010101" => rgb <= "000000";
                when "00011110010110" => rgb <= "000000";
                when "00011110010111" => rgb <= "000000";
                when "00011110011000" => rgb <= "000000";
                when "00011110011001" => rgb <= "000000";
                when "00011110011010" => rgb <= "000000";
                when "00011110011011" => rgb <= "000000";
                when "00011110011100" => rgb <= "000000";
                when "00011110011101" => rgb <= "000000";
                when "00011110011110" => rgb <= "000000";
                when "00011110011111" => rgb <= "000011";
                when "00011110100000" => rgb <= "000011";
                when "00011110100001" => rgb <= "000011";
                when "00011110100010" => rgb <= "000011";
                when "00100000000000" => rgb <= "000000";
                when "00100000000001" => rgb <= "000000";
                when "00100000000010" => rgb <= "000000";
                when "00100000000011" => rgb <= "000000";
                when "00100000000100" => rgb <= "000000";
                when "00100000000101" => rgb <= "000000";
                when "00100000000110" => rgb <= "000000";
                when "00100000000111" => rgb <= "000000";
                when "00100000001000" => rgb <= "000000";
                when "00100000001001" => rgb <= "000000";
                when "00100000001010" => rgb <= "000000";
                when "00100000001011" => rgb <= "000000";
                when "00100000001100" => rgb <= "000000";
                when "00100000001101" => rgb <= "000000";
                when "00100000001110" => rgb <= "000000";
                when "00100000001111" => rgb <= "000000";
                when "00100000010000" => rgb <= "000000";
                when "00100000010001" => rgb <= "000000";
                when "00100000010010" => rgb <= "000000";
                when "00100000010011" => rgb <= "000000";
                when "00100000010100" => rgb <= "000000";
                when "00100000010101" => rgb <= "000000";
                when "00100000010110" => rgb <= "000000";
                when "00100000010111" => rgb <= "000000";
                when "00100000011000" => rgb <= "000000";
                when "00100000011001" => rgb <= "000000";
                when "00100000011010" => rgb <= "000000";
                when "00100000011011" => rgb <= "000000";
                when "00100000011100" => rgb <= "000000";
                when "00100000011101" => rgb <= "000000";
                when "00100000011110" => rgb <= "000000";
                when "00100000011111" => rgb <= "000011";
                when "00100000100000" => rgb <= "000011";
                when "00100000100001" => rgb <= "000011";
                when "00100000100010" => rgb <= "000011";
                when "00100010000000" => rgb <= "000000";
                when "00100010000001" => rgb <= "000000";
                when "00100010000010" => rgb <= "000000";
                when "00100010000011" => rgb <= "000000";
                when "00100010000100" => rgb <= "000000";
                when "00100010000101" => rgb <= "000000";
                when "00100010000110" => rgb <= "000000";
                when "00100010000111" => rgb <= "000000";
                when "00100010001000" => rgb <= "000000";
                when "00100010001001" => rgb <= "000000";
                when "00100010001010" => rgb <= "000000";
                when "00100010001011" => rgb <= "000000";
                when "00100010001100" => rgb <= "000000";
                when "00100010001101" => rgb <= "000000";
                when "00100010001110" => rgb <= "000000";
                when "00100010001111" => rgb <= "000000";
                when "00100010010000" => rgb <= "000000";
                when "00100010010001" => rgb <= "000000";
                when "00100010010010" => rgb <= "000000";
                when "00100010010011" => rgb <= "000000";
                when "00100010010100" => rgb <= "000000";
                when "00100010010101" => rgb <= "000000";
                when "00100010010110" => rgb <= "000000";
                when "00100010010111" => rgb <= "000000";
                when "00100010011000" => rgb <= "000000";
                when "00100010011001" => rgb <= "000000";
                when "00100010011010" => rgb <= "000000";
                when "00100010011011" => rgb <= "000000";
                when "00100010011100" => rgb <= "000000";
                when "00100010011101" => rgb <= "000000";
                when "00100010011110" => rgb <= "000000";
                when "00100010011111" => rgb <= "000011";
                when "00100010100000" => rgb <= "000011";
                when "00100010100001" => rgb <= "000011";
                when "00100010100010" => rgb <= "000011";
                when "00100100000000" => rgb <= "000000";
                when "00100100000001" => rgb <= "000000";
                when "00100100000010" => rgb <= "000000";
                when "00100100000011" => rgb <= "000000";
                when "00100100000100" => rgb <= "000000";
                when "00100100000101" => rgb <= "000000";
                when "00100100000110" => rgb <= "000000";
                when "00100100000111" => rgb <= "000000";
                when "00100100001000" => rgb <= "000000";
                when "00100100001001" => rgb <= "000000";
                when "00100100001010" => rgb <= "000000";
                when "00100100001011" => rgb <= "000000";
                when "00100100001100" => rgb <= "000000";
                when "00100100001101" => rgb <= "000000";
                when "00100100001110" => rgb <= "000000";
                when "00100100001111" => rgb <= "000000";
                when "00100100010000" => rgb <= "000000";
                when "00100100010001" => rgb <= "000000";
                when "00100100010010" => rgb <= "000000";
                when "00100100010011" => rgb <= "000000";
                when "00100100010100" => rgb <= "000000";
                when "00100100010101" => rgb <= "000000";
                when "00100100010110" => rgb <= "000000";
                when "00100100010111" => rgb <= "000000";
                when "00100100011000" => rgb <= "000000";
                when "00100100011001" => rgb <= "000000";
                when "00100100011010" => rgb <= "000000";
                when "00100100011011" => rgb <= "000000";
                when "00100100011100" => rgb <= "000000";
                when "00100100011101" => rgb <= "000000";
                when "00100100011110" => rgb <= "000000";
                when "00100100011111" => rgb <= "000011";
                when "00100100100000" => rgb <= "000011";
                when "00100100100001" => rgb <= "000011";
                when "00100100100010" => rgb <= "000011";
                when "00100110000000" => rgb <= "000000";
                when "00100110000001" => rgb <= "000000";
                when "00100110000010" => rgb <= "000000";
                when "00100110000011" => rgb <= "000000";
                when "00100110000100" => rgb <= "000000";
                when "00100110000101" => rgb <= "000000";
                when "00100110000110" => rgb <= "000000";
                when "00100110000111" => rgb <= "000000";
                when "00100110001000" => rgb <= "000000";
                when "00100110001001" => rgb <= "000000";
                when "00100110001010" => rgb <= "000000";
                when "00100110001011" => rgb <= "000000";
                when "00100110001100" => rgb <= "000000";
                when "00100110001101" => rgb <= "000000";
                when "00100110001110" => rgb <= "000000";
                when "00100110001111" => rgb <= "000000";
                when "00100110010000" => rgb <= "000000";
                when "00100110010001" => rgb <= "000000";
                when "00100110010010" => rgb <= "000000";
                when "00100110010011" => rgb <= "000000";
                when "00100110010100" => rgb <= "000000";
                when "00100110010101" => rgb <= "000000";
                when "00100110010110" => rgb <= "000000";
                when "00100110010111" => rgb <= "000000";
                when "00100110011000" => rgb <= "000000";
                when "00100110011001" => rgb <= "000000";
                when "00100110011010" => rgb <= "000000";
                when "00100110011011" => rgb <= "000000";
                when "00100110011100" => rgb <= "000000";
                when "00100110011101" => rgb <= "000000";
                when "00100110011110" => rgb <= "000000";
                when "00100110011111" => rgb <= "000011";
                when "00100110100000" => rgb <= "000011";
                when "00100110100001" => rgb <= "000011";
                when "00100110100010" => rgb <= "000011";
                when "00101000000000" => rgb <= "000000";
                when "00101000000001" => rgb <= "000000";
                when "00101000000010" => rgb <= "000000";
                when "00101000000011" => rgb <= "000000";
                when "00101000000100" => rgb <= "000000";
                when "00101000000101" => rgb <= "000000";
                when "00101000000110" => rgb <= "000000";
                when "00101000000111" => rgb <= "000000";
                when "00101000001000" => rgb <= "000000";
                when "00101000001001" => rgb <= "000000";
                when "00101000001010" => rgb <= "000000";
                when "00101000001011" => rgb <= "000000";
                when "00101000001100" => rgb <= "000000";
                when "00101000001101" => rgb <= "000000";
                when "00101000001110" => rgb <= "000000";
                when "00101000001111" => rgb <= "000000";
                when "00101000010000" => rgb <= "000000";
                when "00101000010001" => rgb <= "000000";
                when "00101000010010" => rgb <= "000000";
                when "00101000010011" => rgb <= "000000";
                when "00101000010100" => rgb <= "000000";
                when "00101000010101" => rgb <= "000000";
                when "00101000010110" => rgb <= "000000";
                when "00101000010111" => rgb <= "000000";
                when "00101000011000" => rgb <= "000000";
                when "00101000011001" => rgb <= "000000";
                when "00101000011010" => rgb <= "000000";
                when "00101000011011" => rgb <= "000000";
                when "00101000011100" => rgb <= "000000";
                when "00101000011101" => rgb <= "000000";
                when "00101000011110" => rgb <= "000000";
                when "00101000011111" => rgb <= "000011";
                when "00101000100000" => rgb <= "000011";
                when "00101000100001" => rgb <= "000011";
                when "00101000100010" => rgb <= "000011";
                when "00101010000000" => rgb <= "000000";
                when "00101010000001" => rgb <= "000000";
                when "00101010000010" => rgb <= "000000";
                when "00101010000011" => rgb <= "000000";
                when "00101010000100" => rgb <= "000000";
                when "00101010000101" => rgb <= "000000";
                when "00101010000110" => rgb <= "000000";
                when "00101010000111" => rgb <= "000000";
                when "00101010001000" => rgb <= "000000";
                when "00101010001001" => rgb <= "000000";
                when "00101010001010" => rgb <= "000000";
                when "00101010001011" => rgb <= "000000";
                when "00101010001100" => rgb <= "000000";
                when "00101010001101" => rgb <= "000000";
                when "00101010001110" => rgb <= "000000";
                when "00101010001111" => rgb <= "000000";
                when "00101010010000" => rgb <= "000000";
                when "00101010010001" => rgb <= "000000";
                when "00101010010010" => rgb <= "000000";
                when "00101010010011" => rgb <= "000000";
                when "00101010010100" => rgb <= "000000";
                when "00101010010101" => rgb <= "000000";
                when "00101010010110" => rgb <= "000000";
                when "00101010010111" => rgb <= "000000";
                when "00101010011000" => rgb <= "000000";
                when "00101010011001" => rgb <= "000000";
                when "00101010011010" => rgb <= "000000";
                when "00101010011011" => rgb <= "000000";
                when "00101010011100" => rgb <= "000000";
                when "00101010011101" => rgb <= "000000";
                when "00101010011110" => rgb <= "000000";
                when "00101010011111" => rgb <= "000011";
                when "00101010100000" => rgb <= "000011";
                when "00101010100001" => rgb <= "000011";
                when "00101010100010" => rgb <= "000011";
                when "00101100000000" => rgb <= "000000";
                when "00101100000001" => rgb <= "000000";
                when "00101100000010" => rgb <= "000000";
                when "00101100000011" => rgb <= "000000";
                when "00101100000100" => rgb <= "000000";
                when "00101100000101" => rgb <= "000000";
                when "00101100000110" => rgb <= "000000";
                when "00101100000111" => rgb <= "000000";
                when "00101100001000" => rgb <= "000000";
                when "00101100001001" => rgb <= "000000";
                when "00101100001010" => rgb <= "000000";
                when "00101100001011" => rgb <= "000000";
                when "00101100001100" => rgb <= "000000";
                when "00101100001101" => rgb <= "000000";
                when "00101100001110" => rgb <= "000000";
                when "00101100001111" => rgb <= "000000";
                when "00101100010000" => rgb <= "000000";
                when "00101100010001" => rgb <= "000000";
                when "00101100010010" => rgb <= "000000";
                when "00101100010011" => rgb <= "000000";
                when "00101100010100" => rgb <= "000000";
                when "00101100010101" => rgb <= "000000";
                when "00101100010110" => rgb <= "000000";
                when "00101100010111" => rgb <= "000000";
                when "00101100011000" => rgb <= "000000";
                when "00101100011001" => rgb <= "000000";
                when "00101100011010" => rgb <= "000000";
                when "00101100011011" => rgb <= "000000";
                when "00101100011100" => rgb <= "000000";
                when "00101100011101" => rgb <= "000000";
                when "00101100011110" => rgb <= "000000";
                when "00101100011111" => rgb <= "000011";
                when "00101100100000" => rgb <= "000011";
                when "00101100100001" => rgb <= "000011";
                when "00101100100010" => rgb <= "000011";
                when "00101110000000" => rgb <= "000000";
                when "00101110000001" => rgb <= "000000";
                when "00101110000010" => rgb <= "000000";
                when "00101110000011" => rgb <= "000000";
                when "00101110000100" => rgb <= "000000";
                when "00101110000101" => rgb <= "000000";
                when "00101110000110" => rgb <= "000000";
                when "00101110000111" => rgb <= "000000";
                when "00101110001000" => rgb <= "000000";
                when "00101110001001" => rgb <= "000000";
                when "00101110001010" => rgb <= "000000";
                when "00101110001011" => rgb <= "000000";
                when "00101110001100" => rgb <= "000000";
                when "00101110001101" => rgb <= "000000";
                when "00101110001110" => rgb <= "000000";
                when "00101110001111" => rgb <= "000000";
                when "00101110010000" => rgb <= "000000";
                when "00101110010001" => rgb <= "000000";
                when "00101110010010" => rgb <= "000000";
                when "00101110010011" => rgb <= "000000";
                when "00101110010100" => rgb <= "000000";
                when "00101110010101" => rgb <= "000000";
                when "00101110010110" => rgb <= "000000";
                when "00101110010111" => rgb <= "000000";
                when "00101110011000" => rgb <= "000000";
                when "00101110011001" => rgb <= "000000";
                when "00101110011010" => rgb <= "000000";
                when "00101110011011" => rgb <= "000000";
                when "00101110011100" => rgb <= "000000";
                when "00101110011101" => rgb <= "000000";
                when "00101110011110" => rgb <= "000000";
                when "00101110011111" => rgb <= "000011";
                when "00101110100000" => rgb <= "000011";
                when "00101110100001" => rgb <= "000011";
                when "00101110100010" => rgb <= "000011";
                when "00110000000000" => rgb <= "000000";
                when "00110000000001" => rgb <= "000000";
                when "00110000000010" => rgb <= "000000";
                when "00110000000011" => rgb <= "000000";
                when "00110000000100" => rgb <= "000000";
                when "00110000000101" => rgb <= "000000";
                when "00110000000110" => rgb <= "000000";
                when "00110000000111" => rgb <= "000000";
                when "00110000001000" => rgb <= "000000";
                when "00110000001001" => rgb <= "000000";
                when "00110000001010" => rgb <= "000000";
                when "00110000001011" => rgb <= "000000";
                when "00110000001100" => rgb <= "000000";
                when "00110000001101" => rgb <= "000000";
                when "00110000001110" => rgb <= "000000";
                when "00110000001111" => rgb <= "000000";
                when "00110000010000" => rgb <= "000000";
                when "00110000010001" => rgb <= "000000";
                when "00110000010010" => rgb <= "000000";
                when "00110000010011" => rgb <= "000000";
                when "00110000010100" => rgb <= "000000";
                when "00110000010101" => rgb <= "000000";
                when "00110000010110" => rgb <= "000000";
                when "00110000010111" => rgb <= "000000";
                when "00110000011000" => rgb <= "000000";
                when "00110000011001" => rgb <= "000000";
                when "00110000011010" => rgb <= "000000";
                when "00110000011011" => rgb <= "000000";
                when "00110000011100" => rgb <= "000000";
                when "00110000011101" => rgb <= "000000";
                when "00110000011110" => rgb <= "000000";
                when "00110000011111" => rgb <= "000011";
                when "00110000100000" => rgb <= "000011";
                when "00110000100001" => rgb <= "000011";
                when "00110000100010" => rgb <= "000011";
                when "00110010000000" => rgb <= "000000";
                when "00110010000001" => rgb <= "000000";
                when "00110010000010" => rgb <= "000000";
                when "00110010000011" => rgb <= "000000";
                when "00110010000100" => rgb <= "000000";
                when "00110010000101" => rgb <= "000000";
                when "00110010000110" => rgb <= "000000";
                when "00110010000111" => rgb <= "000000";
                when "00110010001000" => rgb <= "000000";
                when "00110010001001" => rgb <= "000000";
                when "00110010001010" => rgb <= "000000";
                when "00110010001011" => rgb <= "000000";
                when "00110010001100" => rgb <= "000000";
                when "00110010001101" => rgb <= "000000";
                when "00110010001110" => rgb <= "000000";
                when "00110010001111" => rgb <= "000000";
                when "00110010010000" => rgb <= "000000";
                when "00110010010001" => rgb <= "000000";
                when "00110010010010" => rgb <= "000000";
                when "00110010010011" => rgb <= "000000";
                when "00110010010100" => rgb <= "000000";
                when "00110010010101" => rgb <= "000000";
                when "00110010010110" => rgb <= "000000";
                when "00110010010111" => rgb <= "000000";
                when "00110010011000" => rgb <= "000000";
                when "00110010011001" => rgb <= "000000";
                when "00110010011010" => rgb <= "000000";
                when "00110010011011" => rgb <= "000000";
                when "00110010011100" => rgb <= "000000";
                when "00110010011101" => rgb <= "000000";
                when "00110010011110" => rgb <= "000000";
                when "00110010011111" => rgb <= "000011";
                when "00110010100000" => rgb <= "000011";
                when "00110010100001" => rgb <= "000011";
                when "00110010100010" => rgb <= "000011";
                when "00110100000000" => rgb <= "000000";
                when "00110100000001" => rgb <= "000000";
                when "00110100000010" => rgb <= "000000";
                when "00110100000011" => rgb <= "000000";
                when "00110100000100" => rgb <= "000000";
                when "00110100000101" => rgb <= "000000";
                when "00110100000110" => rgb <= "000000";
                when "00110100000111" => rgb <= "000000";
                when "00110100001000" => rgb <= "000000";
                when "00110100001001" => rgb <= "000000";
                when "00110100001010" => rgb <= "000000";
                when "00110100001011" => rgb <= "000000";
                when "00110100001100" => rgb <= "000000";
                when "00110100001101" => rgb <= "000000";
                when "00110100001110" => rgb <= "000000";
                when "00110100001111" => rgb <= "000000";
                when "00110100010000" => rgb <= "000000";
                when "00110100010001" => rgb <= "000000";
                when "00110100010010" => rgb <= "000000";
                when "00110100010011" => rgb <= "000000";
                when "00110100010100" => rgb <= "000000";
                when "00110100010101" => rgb <= "000000";
                when "00110100010110" => rgb <= "000000";
                when "00110100010111" => rgb <= "000000";
                when "00110100011000" => rgb <= "000000";
                when "00110100011001" => rgb <= "000000";
                when "00110100011010" => rgb <= "000000";
                when "00110100011011" => rgb <= "000000";
                when "00110100011100" => rgb <= "000000";
                when "00110100011101" => rgb <= "000000";
                when "00110100011110" => rgb <= "000000";
                when "00110100011111" => rgb <= "000011";
                when "00110100100000" => rgb <= "000011";
                when "00110100100001" => rgb <= "000011";
                when "00110100100010" => rgb <= "000011";
                when "00110110000000" => rgb <= "000000";
                when "00110110000001" => rgb <= "000000";
                when "00110110000010" => rgb <= "000000";
                when "00110110000011" => rgb <= "000000";
                when "00110110000100" => rgb <= "000000";
                when "00110110000101" => rgb <= "000000";
                when "00110110000110" => rgb <= "000000";
                when "00110110000111" => rgb <= "000000";
                when "00110110001000" => rgb <= "000000";
                when "00110110001001" => rgb <= "000000";
                when "00110110001010" => rgb <= "000000";
                when "00110110001011" => rgb <= "000000";
                when "00110110001100" => rgb <= "000000";
                when "00110110001101" => rgb <= "000000";
                when "00110110001110" => rgb <= "000000";
                when "00110110001111" => rgb <= "000000";
                when "00110110010000" => rgb <= "000000";
                when "00110110010001" => rgb <= "000000";
                when "00110110010010" => rgb <= "000000";
                when "00110110010011" => rgb <= "000000";
                when "00110110010100" => rgb <= "000000";
                when "00110110010101" => rgb <= "000000";
                when "00110110010110" => rgb <= "000000";
                when "00110110010111" => rgb <= "000000";
                when "00110110011000" => rgb <= "000000";
                when "00110110011001" => rgb <= "000000";
                when "00110110011010" => rgb <= "000000";
                when "00110110011011" => rgb <= "000000";
                when "00110110011100" => rgb <= "000000";
                when "00110110011101" => rgb <= "000000";
                when "00110110011110" => rgb <= "000000";
                when "00110110011111" => rgb <= "000011";
                when "00110110100000" => rgb <= "000011";
                when "00110110100001" => rgb <= "000011";
                when "00110110100010" => rgb <= "000011";
                when "00111000000000" => rgb <= "000000";
                when "00111000000001" => rgb <= "000000";
                when "00111000000010" => rgb <= "000000";
                when "00111000000011" => rgb <= "000000";
                when "00111000000100" => rgb <= "000000";
                when "00111000000101" => rgb <= "000000";
                when "00111000000110" => rgb <= "000000";
                when "00111000000111" => rgb <= "000000";
                when "00111000001000" => rgb <= "000000";
                when "00111000001001" => rgb <= "000000";
                when "00111000001010" => rgb <= "000000";
                when "00111000001011" => rgb <= "000000";
                when "00111000001100" => rgb <= "000000";
                when "00111000001101" => rgb <= "000000";
                when "00111000001110" => rgb <= "000000";
                when "00111000001111" => rgb <= "000000";
                when "00111000010000" => rgb <= "000000";
                when "00111000010001" => rgb <= "000000";
                when "00111000010010" => rgb <= "000000";
                when "00111000010011" => rgb <= "000000";
                when "00111000010100" => rgb <= "000000";
                when "00111000010101" => rgb <= "000000";
                when "00111000010110" => rgb <= "000000";
                when "00111000010111" => rgb <= "000000";
                when "00111000011000" => rgb <= "000000";
                when "00111000011001" => rgb <= "000000";
                when "00111000011010" => rgb <= "000000";
                when "00111000011011" => rgb <= "000000";
                when "00111000011100" => rgb <= "000000";
                when "00111000011101" => rgb <= "000000";
                when "00111000011110" => rgb <= "000000";
                when "00111000011111" => rgb <= "000011";
                when "00111000100000" => rgb <= "000011";
                when "00111000100001" => rgb <= "000011";
                when "00111000100010" => rgb <= "000011";
                when "00111010000000" => rgb <= "000000";
                when "00111010000001" => rgb <= "000000";
                when "00111010000010" => rgb <= "000000";
                when "00111010000011" => rgb <= "000000";
                when "00111010000100" => rgb <= "000000";
                when "00111010000101" => rgb <= "000000";
                when "00111010000110" => rgb <= "000000";
                when "00111010000111" => rgb <= "000000";
                when "00111010001000" => rgb <= "000000";
                when "00111010001001" => rgb <= "000000";
                when "00111010001010" => rgb <= "000000";
                when "00111010001011" => rgb <= "000000";
                when "00111010001100" => rgb <= "000000";
                when "00111010001101" => rgb <= "000000";
                when "00111010001110" => rgb <= "000000";
                when "00111010001111" => rgb <= "000000";
                when "00111010010000" => rgb <= "000000";
                when "00111010010001" => rgb <= "000000";
                when "00111010010010" => rgb <= "000000";
                when "00111010010011" => rgb <= "000000";
                when "00111010010100" => rgb <= "000000";
                when "00111010010101" => rgb <= "000000";
                when "00111010010110" => rgb <= "000000";
                when "00111010010111" => rgb <= "000000";
                when "00111010011000" => rgb <= "000000";
                when "00111010011001" => rgb <= "000000";
                when "00111010011010" => rgb <= "000000";
                when "00111010011011" => rgb <= "000000";
                when "00111010011100" => rgb <= "000000";
                when "00111010011101" => rgb <= "000000";
                when "00111010011110" => rgb <= "000000";
                when "00111010011111" => rgb <= "000011";
                when "00111010100000" => rgb <= "000011";
                when "00111010100001" => rgb <= "000011";
                when "00111010100010" => rgb <= "000011";
                when "00111100000000" => rgb <= "000000";
                when "00111100000001" => rgb <= "000000";
                when "00111100000010" => rgb <= "000000";
                when "00111100000011" => rgb <= "000000";
                when "00111100000100" => rgb <= "000000";
                when "00111100000101" => rgb <= "000000";
                when "00111100000110" => rgb <= "000000";
                when "00111100000111" => rgb <= "000000";
                when "00111100001000" => rgb <= "000000";
                when "00111100001001" => rgb <= "000000";
                when "00111100001010" => rgb <= "000000";
                when "00111100001011" => rgb <= "000000";
                when "00111100001100" => rgb <= "000000";
                when "00111100001101" => rgb <= "000000";
                when "00111100001110" => rgb <= "000000";
                when "00111100001111" => rgb <= "000000";
                when "00111100010000" => rgb <= "000000";
                when "00111100010001" => rgb <= "000000";
                when "00111100010010" => rgb <= "000000";
                when "00111100010011" => rgb <= "000000";
                when "00111100010100" => rgb <= "000000";
                when "00111100010101" => rgb <= "000000";
                when "00111100010110" => rgb <= "000000";
                when "00111100010111" => rgb <= "000000";
                when "00111100011000" => rgb <= "000000";
                when "00111100011001" => rgb <= "000000";
                when "00111100011010" => rgb <= "000000";
                when "00111100011011" => rgb <= "000000";
                when "00111100011100" => rgb <= "000000";
                when "00111100011101" => rgb <= "000000";
                when "00111100011110" => rgb <= "000000";
                when "00111100011111" => rgb <= "000011";
                when "00111100100000" => rgb <= "000011";
                when "00111100100001" => rgb <= "000011";
                when "00111100100010" => rgb <= "000011";
                when "00111110000000" => rgb <= "000000";
                when "00111110000001" => rgb <= "000000";
                when "00111110000010" => rgb <= "000000";
                when "00111110000011" => rgb <= "000000";
                when "00111110000100" => rgb <= "000000";
                when "00111110000101" => rgb <= "000000";
                when "00111110000110" => rgb <= "000000";
                when "00111110000111" => rgb <= "000000";
                when "00111110001000" => rgb <= "000000";
                when "00111110001001" => rgb <= "000000";
                when "00111110001010" => rgb <= "000000";
                when "00111110001011" => rgb <= "000000";
                when "00111110001100" => rgb <= "000000";
                when "00111110001101" => rgb <= "000000";
                when "00111110001110" => rgb <= "000000";
                when "00111110001111" => rgb <= "000000";
                when "00111110010000" => rgb <= "000000";
                when "00111110010001" => rgb <= "000000";
                when "00111110010010" => rgb <= "000000";
                when "00111110010011" => rgb <= "000000";
                when "00111110010100" => rgb <= "000000";
                when "00111110010101" => rgb <= "000000";
                when "00111110010110" => rgb <= "000000";
                when "00111110010111" => rgb <= "000000";
                when "00111110011000" => rgb <= "000000";
                when "00111110011001" => rgb <= "000000";
                when "00111110011010" => rgb <= "000000";
                when "00111110011011" => rgb <= "000000";
                when "00111110011100" => rgb <= "000000";
                when "00111110011101" => rgb <= "000000";
                when "00111110011110" => rgb <= "000000";
                when "00111110011111" => rgb <= "000011";
                when "00111110100000" => rgb <= "000011";
                when "00111110100001" => rgb <= "000011";
                when "00111110100010" => rgb <= "000011";
                when "01000000000000" => rgb <= "000000";
                when "01000000000001" => rgb <= "000000";
                when "01000000000010" => rgb <= "000000";
                when "01000000000011" => rgb <= "000000";
                when "01000000000100" => rgb <= "000000";
                when "01000000000101" => rgb <= "000000";
                when "01000000000110" => rgb <= "000000";
                when "01000000000111" => rgb <= "000000";
                when "01000000001000" => rgb <= "000000";
                when "01000000001001" => rgb <= "000000";
                when "01000000001010" => rgb <= "000000";
                when "01000000001011" => rgb <= "000000";
                when "01000000001100" => rgb <= "000000";
                when "01000000001101" => rgb <= "000000";
                when "01000000001110" => rgb <= "000000";
                when "01000000001111" => rgb <= "000000";
                when "01000000010000" => rgb <= "000000";
                when "01000000010001" => rgb <= "000000";
                when "01000000010010" => rgb <= "000000";
                when "01000000010011" => rgb <= "000000";
                when "01000000010100" => rgb <= "000000";
                when "01000000010101" => rgb <= "000000";
                when "01000000010110" => rgb <= "000000";
                when "01000000010111" => rgb <= "000000";
                when "01000000011000" => rgb <= "000000";
                when "01000000011001" => rgb <= "000000";
                when "01000000011010" => rgb <= "000000";
                when "01000000011011" => rgb <= "000000";
                when "01000000011100" => rgb <= "000000";
                when "01000000011101" => rgb <= "000000";
                when "01000000011110" => rgb <= "000000";
                when "01000000011111" => rgb <= "000011";
                when "01000000100000" => rgb <= "000011";
                when "01000000100001" => rgb <= "000011";
                when "01000000100010" => rgb <= "000011";
                when "01000010000000" => rgb <= "000000";
                when "01000010000001" => rgb <= "000000";
                when "01000010000010" => rgb <= "000000";
                when "01000010000011" => rgb <= "000000";
                when "01000010000100" => rgb <= "000000";
                when "01000010000101" => rgb <= "000000";
                when "01000010000110" => rgb <= "000000";
                when "01000010000111" => rgb <= "000000";
                when "01000010001000" => rgb <= "000000";
                when "01000010001001" => rgb <= "000000";
                when "01000010001010" => rgb <= "000000";
                when "01000010001011" => rgb <= "000000";
                when "01000010001100" => rgb <= "000000";
                when "01000010001101" => rgb <= "000000";
                when "01000010001110" => rgb <= "000000";
                when "01000010001111" => rgb <= "000000";
                when "01000010010000" => rgb <= "000000";
                when "01000010010001" => rgb <= "000000";
                when "01000010010010" => rgb <= "000000";
                when "01000010010011" => rgb <= "000000";
                when "01000010010100" => rgb <= "000000";
                when "01000010010101" => rgb <= "000000";
                when "01000010010110" => rgb <= "000000";
                when "01000010010111" => rgb <= "000000";
                when "01000010011000" => rgb <= "000000";
                when "01000010011001" => rgb <= "000000";
                when "01000010011010" => rgb <= "000000";
                when "01000010011011" => rgb <= "000000";
                when "01000010011100" => rgb <= "000000";
                when "01000010011101" => rgb <= "000000";
                when "01000010011110" => rgb <= "000000";
                when "01000010011111" => rgb <= "000011";
                when "01000010100000" => rgb <= "000011";
                when "01000010100001" => rgb <= "000011";
                when "01000010100010" => rgb <= "000011";
                when "01000100000000" => rgb <= "000000";
                when "01000100000001" => rgb <= "000000";
                when "01000100000010" => rgb <= "000000";
                when "01000100000011" => rgb <= "000000";
                when "01000100000100" => rgb <= "000000";
                when "01000100000101" => rgb <= "000000";
                when "01000100000110" => rgb <= "000000";
                when "01000100000111" => rgb <= "000000";
                when "01000100001000" => rgb <= "000000";
                when "01000100001001" => rgb <= "000000";
                when "01000100001010" => rgb <= "000000";
                when "01000100001011" => rgb <= "000000";
                when "01000100001100" => rgb <= "000000";
                when "01000100001101" => rgb <= "000000";
                when "01000100001110" => rgb <= "000000";
                when "01000100001111" => rgb <= "000000";
                when "01000100010000" => rgb <= "000000";
                when "01000100010001" => rgb <= "000000";
                when "01000100010010" => rgb <= "000000";
                when "01000100010011" => rgb <= "000000";
                when "01000100010100" => rgb <= "000000";
                when "01000100010101" => rgb <= "000000";
                when "01000100010110" => rgb <= "000000";
                when "01000100010111" => rgb <= "000000";
                when "01000100011000" => rgb <= "000000";
                when "01000100011001" => rgb <= "000000";
                when "01000100011010" => rgb <= "000000";
                when "01000100011011" => rgb <= "000000";
                when "01000100011100" => rgb <= "000000";
                when "01000100011101" => rgb <= "000000";
                when "01000100011110" => rgb <= "000000";
                when "01000100011111" => rgb <= "000011";
                when "01000100100000" => rgb <= "000011";
                when "01000100100001" => rgb <= "000011";
                when "01000100100010" => rgb <= "000011";
                when "01000110000000" => rgb <= "000000";
                when "01000110000001" => rgb <= "000000";
                when "01000110000010" => rgb <= "000000";
                when "01000110000011" => rgb <= "000000";
                when "01000110000100" => rgb <= "000000";
                when "01000110000101" => rgb <= "000000";
                when "01000110000110" => rgb <= "000000";
                when "01000110000111" => rgb <= "000000";
                when "01000110001000" => rgb <= "000000";
                when "01000110001001" => rgb <= "000000";
                when "01000110001010" => rgb <= "000000";
                when "01000110001011" => rgb <= "000000";
                when "01000110001100" => rgb <= "000000";
                when "01000110001101" => rgb <= "000000";
                when "01000110001110" => rgb <= "000000";
                when "01000110001111" => rgb <= "000000";
                when "01000110010000" => rgb <= "000000";
                when "01000110010001" => rgb <= "000000";
                when "01000110010010" => rgb <= "000000";
                when "01000110010011" => rgb <= "000000";
                when "01000110010100" => rgb <= "000000";
                when "01000110010101" => rgb <= "000000";
                when "01000110010110" => rgb <= "000000";
                when "01000110010111" => rgb <= "000000";
                when "01000110011000" => rgb <= "000000";
                when "01000110011001" => rgb <= "000000";
                when "01000110011010" => rgb <= "000000";
                when "01000110011011" => rgb <= "000000";
                when "01000110011100" => rgb <= "000000";
                when "01000110011101" => rgb <= "000000";
                when "01000110011110" => rgb <= "000000";
                when "01000110011111" => rgb <= "000011";
                when "01000110100000" => rgb <= "000011";
                when "01000110100001" => rgb <= "000011";
                when "01000110100010" => rgb <= "000011";
                when "01001000000000" => rgb <= "000000";
                when "01001000000001" => rgb <= "000000";
                when "01001000000010" => rgb <= "000000";
                when "01001000000011" => rgb <= "000000";
                when "01001000000100" => rgb <= "000000";
                when "01001000000101" => rgb <= "000000";
                when "01001000000110" => rgb <= "000000";
                when "01001000000111" => rgb <= "000000";
                when "01001000001000" => rgb <= "000000";
                when "01001000001001" => rgb <= "000000";
                when "01001000001010" => rgb <= "000000";
                when "01001000001011" => rgb <= "000000";
                when "01001000001100" => rgb <= "000000";
                when "01001000001101" => rgb <= "000000";
                when "01001000001110" => rgb <= "000000";
                when "01001000001111" => rgb <= "000000";
                when "01001000010000" => rgb <= "000000";
                when "01001000010001" => rgb <= "000000";
                when "01001000010010" => rgb <= "000000";
                when "01001000010011" => rgb <= "000000";
                when "01001000010100" => rgb <= "000000";
                when "01001000010101" => rgb <= "000000";
                when "01001000010110" => rgb <= "000000";
                when "01001000010111" => rgb <= "000000";
                when "01001000011000" => rgb <= "000000";
                when "01001000011001" => rgb <= "000000";
                when "01001000011010" => rgb <= "000000";
                when "01001000011011" => rgb <= "000000";
                when "01001000011100" => rgb <= "000000";
                when "01001000011101" => rgb <= "000000";
                when "01001000011110" => rgb <= "000000";
                when "01001000011111" => rgb <= "000011";
                when "01001000100000" => rgb <= "000011";
                when "01001000100001" => rgb <= "000011";
                when "01001000100010" => rgb <= "000011";
                when "01001010000000" => rgb <= "000000";
                when "01001010000001" => rgb <= "000000";
                when "01001010000010" => rgb <= "000000";
                when "01001010000011" => rgb <= "000000";
                when "01001010000100" => rgb <= "000000";
                when "01001010000101" => rgb <= "000000";
                when "01001010000110" => rgb <= "000000";
                when "01001010000111" => rgb <= "000000";
                when "01001010001000" => rgb <= "000000";
                when "01001010001001" => rgb <= "000000";
                when "01001010001010" => rgb <= "000000";
                when "01001010001011" => rgb <= "000000";
                when "01001010001100" => rgb <= "000000";
                when "01001010001101" => rgb <= "000000";
                when "01001010001110" => rgb <= "000000";
                when "01001010001111" => rgb <= "000000";
                when "01001010010000" => rgb <= "000000";
                when "01001010010001" => rgb <= "000000";
                when "01001010010010" => rgb <= "000000";
                when "01001010010011" => rgb <= "000000";
                when "01001010010100" => rgb <= "000000";
                when "01001010010101" => rgb <= "000000";
                when "01001010010110" => rgb <= "000000";
                when "01001010010111" => rgb <= "000000";
                when "01001010011000" => rgb <= "000000";
                when "01001010011001" => rgb <= "000000";
                when "01001010011010" => rgb <= "000000";
                when "01001010011011" => rgb <= "000000";
                when "01001010011100" => rgb <= "000000";
                when "01001010011101" => rgb <= "000000";
                when "01001010011110" => rgb <= "000000";
                when "01001010011111" => rgb <= "000011";
                when "01001010100000" => rgb <= "000011";
                when "01001010100001" => rgb <= "000011";
                when "01001010100010" => rgb <= "000011";
                when "01001100000000" => rgb <= "000000";
                when "01001100000001" => rgb <= "000000";
                when "01001100000010" => rgb <= "000000";
                when "01001100000011" => rgb <= "000000";
                when "01001100000100" => rgb <= "000000";
                when "01001100000101" => rgb <= "000000";
                when "01001100000110" => rgb <= "000000";
                when "01001100000111" => rgb <= "000000";
                when "01001100001000" => rgb <= "000000";
                when "01001100001001" => rgb <= "000000";
                when "01001100001010" => rgb <= "000000";
                when "01001100001011" => rgb <= "000000";
                when "01001100001100" => rgb <= "000000";
                when "01001100001101" => rgb <= "000000";
                when "01001100001110" => rgb <= "000000";
                when "01001100001111" => rgb <= "000000";
                when "01001100010000" => rgb <= "000000";
                when "01001100010001" => rgb <= "000000";
                when "01001100010010" => rgb <= "000000";
                when "01001100010011" => rgb <= "000000";
                when "01001100010100" => rgb <= "000000";
                when "01001100010101" => rgb <= "000000";
                when "01001100010110" => rgb <= "000000";
                when "01001100010111" => rgb <= "000000";
                when "01001100011000" => rgb <= "000000";
                when "01001100011001" => rgb <= "000000";
                when "01001100011010" => rgb <= "000000";
                when "01001100011011" => rgb <= "000000";
                when "01001100011100" => rgb <= "000000";
                when "01001100011101" => rgb <= "000000";
                when "01001100011110" => rgb <= "000000";
                when "01001100011111" => rgb <= "000011";
                when "01001100100000" => rgb <= "000011";
                when "01001100100001" => rgb <= "000011";
                when "01001100100010" => rgb <= "000011";
                when "01001110000000" => rgb <= "000000";
                when "01001110000001" => rgb <= "000000";
                when "01001110000010" => rgb <= "000000";
                when "01001110000011" => rgb <= "000000";
                when "01001110000100" => rgb <= "000000";
                when "01001110000101" => rgb <= "000000";
                when "01001110000110" => rgb <= "000000";
                when "01001110000111" => rgb <= "000000";
                when "01001110001000" => rgb <= "000000";
                when "01001110001001" => rgb <= "000000";
                when "01001110001010" => rgb <= "000000";
                when "01001110001011" => rgb <= "000000";
                when "01001110001100" => rgb <= "000000";
                when "01001110001101" => rgb <= "000000";
                when "01001110001110" => rgb <= "000000";
                when "01001110001111" => rgb <= "000000";
                when "01001110010000" => rgb <= "000000";
                when "01001110010001" => rgb <= "000000";
                when "01001110010010" => rgb <= "000000";
                when "01001110010011" => rgb <= "000000";
                when "01001110010100" => rgb <= "000000";
                when "01001110010101" => rgb <= "000000";
                when "01001110010110" => rgb <= "000000";
                when "01001110010111" => rgb <= "000000";
                when "01001110011000" => rgb <= "000000";
                when "01001110011001" => rgb <= "000000";
                when "01001110011010" => rgb <= "000000";
                when "01001110011011" => rgb <= "000000";
                when "01001110011100" => rgb <= "000000";
                when "01001110011101" => rgb <= "000000";
                when "01001110011110" => rgb <= "000000";
                when "01001110011111" => rgb <= "000011";
                when "01001110100000" => rgb <= "000011";
                when "01001110100001" => rgb <= "000011";
                when "01001110100010" => rgb <= "000011";
                when "01010000000000" => rgb <= "000000";
                when "01010000000001" => rgb <= "000000";
                when "01010000000010" => rgb <= "000000";
                when "01010000000011" => rgb <= "000000";
                when "01010000000100" => rgb <= "000000";
                when "01010000000101" => rgb <= "000000";
                when "01010000000110" => rgb <= "000000";
                when "01010000000111" => rgb <= "000000";
                when "01010000001000" => rgb <= "000000";
                when "01010000001001" => rgb <= "000000";
                when "01010000001010" => rgb <= "000000";
                when "01010000001011" => rgb <= "000000";
                when "01010000001100" => rgb <= "000000";
                when "01010000001101" => rgb <= "000000";
                when "01010000001110" => rgb <= "000000";
                when "01010000001111" => rgb <= "000000";
                when "01010000010000" => rgb <= "000000";
                when "01010000010001" => rgb <= "000000";
                when "01010000010010" => rgb <= "000000";
                when "01010000010011" => rgb <= "000000";
                when "01010000010100" => rgb <= "000000";
                when "01010000010101" => rgb <= "000000";
                when "01010000010110" => rgb <= "000000";
                when "01010000010111" => rgb <= "000000";
                when "01010000011000" => rgb <= "000000";
                when "01010000011001" => rgb <= "000000";
                when "01010000011010" => rgb <= "000000";
                when "01010000011011" => rgb <= "000000";
                when "01010000011100" => rgb <= "000000";
                when "01010000011101" => rgb <= "000000";
                when "01010000011110" => rgb <= "000000";
                when "01010000011111" => rgb <= "000011";
                when "01010000100000" => rgb <= "000011";
                when "01010000100001" => rgb <= "000011";
                when "01010000100010" => rgb <= "000011";
                when "01010010000000" => rgb <= "000000";
                when "01010010000001" => rgb <= "000000";
                when "01010010000010" => rgb <= "000000";
                when "01010010000011" => rgb <= "000000";
                when "01010010000100" => rgb <= "000000";
                when "01010010000101" => rgb <= "000000";
                when "01010010000110" => rgb <= "000000";
                when "01010010000111" => rgb <= "000000";
                when "01010010001000" => rgb <= "000000";
                when "01010010001001" => rgb <= "000000";
                when "01010010001010" => rgb <= "000000";
                when "01010010001011" => rgb <= "000000";
                when "01010010001100" => rgb <= "000000";
                when "01010010001101" => rgb <= "000000";
                when "01010010001110" => rgb <= "000000";
                when "01010010001111" => rgb <= "000000";
                when "01010010010000" => rgb <= "000000";
                when "01010010010001" => rgb <= "000000";
                when "01010010010010" => rgb <= "000000";
                when "01010010010011" => rgb <= "000000";
                when "01010010010100" => rgb <= "000000";
                when "01010010010101" => rgb <= "000000";
                when "01010010010110" => rgb <= "000000";
                when "01010010010111" => rgb <= "000000";
                when "01010010011000" => rgb <= "000000";
                when "01010010011001" => rgb <= "000000";
                when "01010010011010" => rgb <= "000000";
                when "01010010011011" => rgb <= "000000";
                when "01010010011100" => rgb <= "000000";
                when "01010010011101" => rgb <= "000000";
                when "01010010011110" => rgb <= "000000";
                when "01010010011111" => rgb <= "000011";
                when "01010010100000" => rgb <= "000011";
                when "01010010100001" => rgb <= "000011";
                when "01010010100010" => rgb <= "000011";
                when "01010100000000" => rgb <= "000000";
                when "01010100000001" => rgb <= "000000";
                when "01010100000010" => rgb <= "000000";
                when "01010100000011" => rgb <= "000000";
                when "01010100000100" => rgb <= "000000";
                when "01010100000101" => rgb <= "000000";
                when "01010100000110" => rgb <= "000000";
                when "01010100000111" => rgb <= "000000";
                when "01010100001000" => rgb <= "000000";
                when "01010100001001" => rgb <= "000000";
                when "01010100001010" => rgb <= "000000";
                when "01010100001011" => rgb <= "000000";
                when "01010100001100" => rgb <= "000000";
                when "01010100001101" => rgb <= "000000";
                when "01010100001110" => rgb <= "000000";
                when "01010100001111" => rgb <= "000000";
                when "01010100010000" => rgb <= "000000";
                when "01010100010001" => rgb <= "000000";
                when "01010100010010" => rgb <= "000000";
                when "01010100010011" => rgb <= "000000";
                when "01010100010100" => rgb <= "000000";
                when "01010100010101" => rgb <= "000000";
                when "01010100010110" => rgb <= "000000";
                when "01010100010111" => rgb <= "000000";
                when "01010100011000" => rgb <= "000000";
                when "01010100011001" => rgb <= "000000";
                when "01010100011010" => rgb <= "000000";
                when "01010100011011" => rgb <= "000000";
                when "01010100011100" => rgb <= "000000";
                when "01010100011101" => rgb <= "000000";
                when "01010100011110" => rgb <= "000000";
                when "01010100011111" => rgb <= "000011";
                when "01010100100000" => rgb <= "000011";
                when "01010100100001" => rgb <= "000011";
                when "01010100100010" => rgb <= "000011";
                when "01010110000000" => rgb <= "000000";
                when "01010110000001" => rgb <= "000000";
                when "01010110000010" => rgb <= "000000";
                when "01010110000011" => rgb <= "000000";
                when "01010110000100" => rgb <= "000000";
                when "01010110000101" => rgb <= "000000";
                when "01010110000110" => rgb <= "000000";
                when "01010110000111" => rgb <= "000000";
                when "01010110001000" => rgb <= "000000";
                when "01010110001001" => rgb <= "000000";
                when "01010110001010" => rgb <= "000000";
                when "01010110001011" => rgb <= "000000";
                when "01010110001100" => rgb <= "000000";
                when "01010110001101" => rgb <= "000000";
                when "01010110001110" => rgb <= "000000";
                when "01010110001111" => rgb <= "000000";
                when "01010110010000" => rgb <= "000000";
                when "01010110010001" => rgb <= "000000";
                when "01010110010010" => rgb <= "000000";
                when "01010110010011" => rgb <= "000000";
                when "01010110010100" => rgb <= "000000";
                when "01010110010101" => rgb <= "000000";
                when "01010110010110" => rgb <= "000000";
                when "01010110010111" => rgb <= "000000";
                when "01010110011000" => rgb <= "000000";
                when "01010110011001" => rgb <= "000000";
                when "01010110011010" => rgb <= "000000";
                when "01010110011011" => rgb <= "000000";
                when "01010110011100" => rgb <= "000000";
                when "01010110011101" => rgb <= "000000";
                when "01010110011110" => rgb <= "000000";
                when "01010110011111" => rgb <= "000011";
                when "01010110100000" => rgb <= "000011";
                when "01010110100001" => rgb <= "000011";
                when "01010110100010" => rgb <= "000011";
                when "01011000000000" => rgb <= "000000";
                when "01011000000001" => rgb <= "000000";
                when "01011000000010" => rgb <= "000000";
                when "01011000000011" => rgb <= "000000";
                when "01011000000100" => rgb <= "000000";
                when "01011000000101" => rgb <= "000000";
                when "01011000000110" => rgb <= "000000";
                when "01011000000111" => rgb <= "000000";
                when "01011000001000" => rgb <= "000000";
                when "01011000001001" => rgb <= "000000";
                when "01011000001010" => rgb <= "000000";
                when "01011000001011" => rgb <= "000000";
                when "01011000001100" => rgb <= "000000";
                when "01011000001101" => rgb <= "000000";
                when "01011000001110" => rgb <= "000000";
                when "01011000001111" => rgb <= "000000";
                when "01011000010000" => rgb <= "000000";
                when "01011000010001" => rgb <= "000000";
                when "01011000010010" => rgb <= "000000";
                when "01011000010011" => rgb <= "000000";
                when "01011000010100" => rgb <= "000000";
                when "01011000010101" => rgb <= "000000";
                when "01011000010110" => rgb <= "000000";
                when "01011000010111" => rgb <= "000000";
                when "01011000011000" => rgb <= "000000";
                when "01011000011001" => rgb <= "000000";
                when "01011000011010" => rgb <= "000000";
                when "01011000011011" => rgb <= "000000";
                when "01011000011100" => rgb <= "000000";
                when "01011000011101" => rgb <= "000000";
                when "01011000011110" => rgb <= "000000";
                when "01011000011111" => rgb <= "000011";
                when "01011000100000" => rgb <= "000011";
                when "01011000100001" => rgb <= "000011";
                when "01011000100010" => rgb <= "000011";
                when "01011010000000" => rgb <= "000000";
                when "01011010000001" => rgb <= "000000";
                when "01011010000010" => rgb <= "000000";
                when "01011010000011" => rgb <= "000000";
                when "01011010000100" => rgb <= "000000";
                when "01011010000101" => rgb <= "000000";
                when "01011010000110" => rgb <= "000000";
                when "01011010000111" => rgb <= "000000";
                when "01011010001000" => rgb <= "000000";
                when "01011010001001" => rgb <= "000000";
                when "01011010001010" => rgb <= "000000";
                when "01011010001011" => rgb <= "000000";
                when "01011010001100" => rgb <= "000000";
                when "01011010001101" => rgb <= "000000";
                when "01011010001110" => rgb <= "000000";
                when "01011010001111" => rgb <= "000000";
                when "01011010010000" => rgb <= "000000";
                when "01011010010001" => rgb <= "000000";
                when "01011010010010" => rgb <= "000000";
                when "01011010010011" => rgb <= "000000";
                when "01011010010100" => rgb <= "000000";
                when "01011010010101" => rgb <= "000000";
                when "01011010010110" => rgb <= "000000";
                when "01011010010111" => rgb <= "000000";
                when "01011010011000" => rgb <= "000000";
                when "01011010011001" => rgb <= "000000";
                when "01011010011010" => rgb <= "000000";
                when "01011010011011" => rgb <= "000000";
                when "01011010011100" => rgb <= "000000";
                when "01011010011101" => rgb <= "000000";
                when "01011010011110" => rgb <= "000000";
                when "01011010011111" => rgb <= "000011";
                when "01011010100000" => rgb <= "000011";
                when "01011010100001" => rgb <= "000011";
                when "01011010100010" => rgb <= "000011";
                when "01011100000000" => rgb <= "000000";
                when "01011100000001" => rgb <= "000000";
                when "01011100000010" => rgb <= "000000";
                when "01011100000011" => rgb <= "000000";
                when "01011100000100" => rgb <= "000000";
                when "01011100000101" => rgb <= "000000";
                when "01011100000110" => rgb <= "000000";
                when "01011100000111" => rgb <= "000000";
                when "01011100001000" => rgb <= "000000";
                when "01011100001001" => rgb <= "000000";
                when "01011100001010" => rgb <= "000000";
                when "01011100001011" => rgb <= "000000";
                when "01011100001100" => rgb <= "000000";
                when "01011100001101" => rgb <= "000000";
                when "01011100001110" => rgb <= "000000";
                when "01011100001111" => rgb <= "000000";
                when "01011100010000" => rgb <= "000000";
                when "01011100010001" => rgb <= "000000";
                when "01011100010010" => rgb <= "000000";
                when "01011100010011" => rgb <= "000000";
                when "01011100010100" => rgb <= "000000";
                when "01011100010101" => rgb <= "000000";
                when "01011100010110" => rgb <= "000000";
                when "01011100010111" => rgb <= "000000";
                when "01011100011000" => rgb <= "000000";
                when "01011100011001" => rgb <= "000000";
                when "01011100011010" => rgb <= "000000";
                when "01011100011011" => rgb <= "000000";
                when "01011100011100" => rgb <= "000000";
                when "01011100011101" => rgb <= "000000";
                when "01011100011110" => rgb <= "000000";
                when "01011100011111" => rgb <= "000011";
                when "01011100100000" => rgb <= "000011";
                when "01011100100001" => rgb <= "000011";
                when "01011100100010" => rgb <= "000011";
                when "01011110000000" => rgb <= "000000";
                when "01011110000001" => rgb <= "000000";
                when "01011110000010" => rgb <= "000000";
                when "01011110000011" => rgb <= "000000";
                when "01011110000100" => rgb <= "000000";
                when "01011110000101" => rgb <= "000000";
                when "01011110000110" => rgb <= "000000";
                when "01011110000111" => rgb <= "000000";
                when "01011110001000" => rgb <= "000000";
                when "01011110001001" => rgb <= "000000";
                when "01011110001010" => rgb <= "000000";
                when "01011110001011" => rgb <= "000000";
                when "01011110001100" => rgb <= "000000";
                when "01011110001101" => rgb <= "000000";
                when "01011110001110" => rgb <= "000000";
                when "01011110001111" => rgb <= "000000";
                when "01011110010000" => rgb <= "000000";
                when "01011110010001" => rgb <= "000000";
                when "01011110010010" => rgb <= "000000";
                when "01011110010011" => rgb <= "000000";
                when "01011110010100" => rgb <= "000000";
                when "01011110010101" => rgb <= "000000";
                when "01011110010110" => rgb <= "000000";
                when "01011110010111" => rgb <= "000000";
                when "01011110011000" => rgb <= "000000";
                when "01011110011001" => rgb <= "000000";
                when "01011110011010" => rgb <= "000000";
                when "01011110011011" => rgb <= "000000";
                when "01011110011100" => rgb <= "000000";
                when "01011110011101" => rgb <= "000000";
                when "01011110011110" => rgb <= "000000";
                when "01011110011111" => rgb <= "000011";
                when "01011110100000" => rgb <= "000011";
                when "01011110100001" => rgb <= "000011";
                when "01011110100010" => rgb <= "000011";
                when "01100000000000" => rgb <= "000000";
                when "01100000000001" => rgb <= "000000";
                when "01100000000010" => rgb <= "000000";
                when "01100000000011" => rgb <= "000000";
                when "01100000000100" => rgb <= "000000";
                when "01100000000101" => rgb <= "000000";
                when "01100000000110" => rgb <= "000000";
                when "01100000000111" => rgb <= "000000";
                when "01100000001000" => rgb <= "000000";
                when "01100000001001" => rgb <= "000000";
                when "01100000001010" => rgb <= "000000";
                when "01100000001011" => rgb <= "000000";
                when "01100000001100" => rgb <= "000000";
                when "01100000001101" => rgb <= "000000";
                when "01100000001110" => rgb <= "000000";
                when "01100000001111" => rgb <= "000000";
                when "01100000010000" => rgb <= "000000";
                when "01100000010001" => rgb <= "000000";
                when "01100000010010" => rgb <= "000000";
                when "01100000010011" => rgb <= "000000";
                when "01100000010100" => rgb <= "000000";
                when "01100000010101" => rgb <= "000000";
                when "01100000010110" => rgb <= "000000";
                when "01100000010111" => rgb <= "000000";
                when "01100000011000" => rgb <= "000000";
                when "01100000011001" => rgb <= "000000";
                when "01100000011010" => rgb <= "000000";
                when "01100000011011" => rgb <= "000000";
                when "01100000011100" => rgb <= "000000";
                when "01100000011101" => rgb <= "000000";
                when "01100000011110" => rgb <= "000000";
                when "01100000011111" => rgb <= "000011";
                when "01100000100000" => rgb <= "000011";
                when "01100000100001" => rgb <= "000011";
                when "01100000100010" => rgb <= "000011";
                when "01100010000000" => rgb <= "000000";
                when "01100010000001" => rgb <= "000000";
                when "01100010000010" => rgb <= "000000";
                when "01100010000011" => rgb <= "000000";
                when "01100010000100" => rgb <= "000000";
                when "01100010000101" => rgb <= "000000";
                when "01100010000110" => rgb <= "000000";
                when "01100010000111" => rgb <= "000000";
                when "01100010001000" => rgb <= "000000";
                when "01100010001001" => rgb <= "000000";
                when "01100010001010" => rgb <= "000000";
                when "01100010001011" => rgb <= "000000";
                when "01100010001100" => rgb <= "000000";
                when "01100010001101" => rgb <= "000000";
                when "01100010001110" => rgb <= "000000";
                when "01100010001111" => rgb <= "000000";
                when "01100010010000" => rgb <= "000000";
                when "01100010010001" => rgb <= "000000";
                when "01100010010010" => rgb <= "000000";
                when "01100010010011" => rgb <= "000000";
                when "01100010010100" => rgb <= "000000";
                when "01100010010101" => rgb <= "000000";
                when "01100010010110" => rgb <= "000000";
                when "01100010010111" => rgb <= "000000";
                when "01100010011000" => rgb <= "000000";
                when "01100010011001" => rgb <= "000000";
                when "01100010011010" => rgb <= "000000";
                when "01100010011011" => rgb <= "000000";
                when "01100010011100" => rgb <= "000000";
                when "01100010011101" => rgb <= "000000";
                when "01100010011110" => rgb <= "000000";
                when "01100010011111" => rgb <= "000011";
                when "01100010100000" => rgb <= "000011";
                when "01100010100001" => rgb <= "000011";
                when "01100010100010" => rgb <= "000011";
                when "01100100000000" => rgb <= "000000";
                when "01100100000001" => rgb <= "000000";
                when "01100100000010" => rgb <= "000000";
                when "01100100000011" => rgb <= "000000";
                when "01100100000100" => rgb <= "000000";
                when "01100100000101" => rgb <= "000000";
                when "01100100000110" => rgb <= "000000";
                when "01100100000111" => rgb <= "000000";
                when "01100100001000" => rgb <= "000000";
                when "01100100001001" => rgb <= "000000";
                when "01100100001010" => rgb <= "000000";
                when "01100100001011" => rgb <= "000000";
                when "01100100001100" => rgb <= "000000";
                when "01100100001101" => rgb <= "000000";
                when "01100100001110" => rgb <= "000000";
                when "01100100001111" => rgb <= "000000";
                when "01100100010000" => rgb <= "000000";
                when "01100100010001" => rgb <= "000000";
                when "01100100010010" => rgb <= "000000";
                when "01100100010011" => rgb <= "000000";
                when "01100100010100" => rgb <= "000000";
                when "01100100010101" => rgb <= "000000";
                when "01100100010110" => rgb <= "000000";
                when "01100100010111" => rgb <= "000000";
                when "01100100011000" => rgb <= "000000";
                when "01100100011001" => rgb <= "000000";
                when "01100100011010" => rgb <= "000000";
                when "01100100011011" => rgb <= "000000";
                when "01100100011100" => rgb <= "000000";
                when "01100100011101" => rgb <= "000000";
                when "01100100011110" => rgb <= "000000";
                when "01100100011111" => rgb <= "000011";
                when "01100100100000" => rgb <= "000011";
                when "01100100100001" => rgb <= "000011";
                when "01100100100010" => rgb <= "000011";
                when "01100110000000" => rgb <= "000000";
                when "01100110000001" => rgb <= "000000";
                when "01100110000010" => rgb <= "000000";
                when "01100110000011" => rgb <= "000000";
                when "01100110000100" => rgb <= "000000";
                when "01100110000101" => rgb <= "000000";
                when "01100110000110" => rgb <= "000000";
                when "01100110000111" => rgb <= "000000";
                when "01100110001000" => rgb <= "000000";
                when "01100110001001" => rgb <= "000000";
                when "01100110001010" => rgb <= "000000";
                when "01100110001011" => rgb <= "000000";
                when "01100110001100" => rgb <= "000000";
                when "01100110001101" => rgb <= "000000";
                when "01100110001110" => rgb <= "000000";
                when "01100110001111" => rgb <= "000000";
                when "01100110010000" => rgb <= "000000";
                when "01100110010001" => rgb <= "000000";
                when "01100110010010" => rgb <= "000000";
                when "01100110010011" => rgb <= "000000";
                when "01100110010100" => rgb <= "000000";
                when "01100110010101" => rgb <= "000000";
                when "01100110010110" => rgb <= "000000";
                when "01100110010111" => rgb <= "000000";
                when "01100110011000" => rgb <= "000000";
                when "01100110011001" => rgb <= "000000";
                when "01100110011010" => rgb <= "000000";
                when "01100110011011" => rgb <= "000000";
                when "01100110011100" => rgb <= "000000";
                when "01100110011101" => rgb <= "000000";
                when "01100110011110" => rgb <= "000000";
                when "01100110011111" => rgb <= "000011";
                when "01100110100000" => rgb <= "000011";
                when "01100110100001" => rgb <= "000011";
                when "01100110100010" => rgb <= "000011";
                when "01101000000000" => rgb <= "000000";
                when "01101000000001" => rgb <= "000000";
                when "01101000000010" => rgb <= "000000";
                when "01101000000011" => rgb <= "000000";
                when "01101000000100" => rgb <= "000000";
                when "01101000000101" => rgb <= "000000";
                when "01101000000110" => rgb <= "000000";
                when "01101000000111" => rgb <= "000000";
                when "01101000001000" => rgb <= "000000";
                when "01101000001001" => rgb <= "000000";
                when "01101000001010" => rgb <= "000000";
                when "01101000001011" => rgb <= "000000";
                when "01101000001100" => rgb <= "000000";
                when "01101000001101" => rgb <= "000000";
                when "01101000001110" => rgb <= "000000";
                when "01101000001111" => rgb <= "000000";
                when "01101000010000" => rgb <= "000000";
                when "01101000010001" => rgb <= "000000";
                when "01101000010010" => rgb <= "000000";
                when "01101000010011" => rgb <= "000000";
                when "01101000010100" => rgb <= "000000";
                when "01101000010101" => rgb <= "000000";
                when "01101000010110" => rgb <= "000000";
                when "01101000010111" => rgb <= "000000";
                when "01101000011000" => rgb <= "000000";
                when "01101000011001" => rgb <= "000000";
                when "01101000011010" => rgb <= "000000";
                when "01101000011011" => rgb <= "000000";
                when "01101000011100" => rgb <= "000000";
                when "01101000011101" => rgb <= "000000";
                when "01101000011110" => rgb <= "000000";
                when "01101000011111" => rgb <= "000011";
                when "01101000100000" => rgb <= "000011";
                when "01101000100001" => rgb <= "000011";
                when "01101000100010" => rgb <= "000011";
                when "01101010000000" => rgb <= "000000";
                when "01101010000001" => rgb <= "000000";
                when "01101010000010" => rgb <= "000000";
                when "01101010000011" => rgb <= "000000";
                when "01101010000100" => rgb <= "000000";
                when "01101010000101" => rgb <= "000000";
                when "01101010000110" => rgb <= "000000";
                when "01101010000111" => rgb <= "000000";
                when "01101010001000" => rgb <= "000000";
                when "01101010001001" => rgb <= "000000";
                when "01101010001010" => rgb <= "000000";
                when "01101010001011" => rgb <= "000000";
                when "01101010001100" => rgb <= "000000";
                when "01101010001101" => rgb <= "000000";
                when "01101010001110" => rgb <= "000000";
                when "01101010001111" => rgb <= "000000";
                when "01101010010000" => rgb <= "000000";
                when "01101010010001" => rgb <= "000000";
                when "01101010010010" => rgb <= "000000";
                when "01101010010011" => rgb <= "000000";
                when "01101010010100" => rgb <= "000000";
                when "01101010010101" => rgb <= "000000";
                when "01101010010110" => rgb <= "000000";
                when "01101010010111" => rgb <= "000000";
                when "01101010011000" => rgb <= "000000";
                when "01101010011001" => rgb <= "000000";
                when "01101010011010" => rgb <= "000000";
                when "01101010011011" => rgb <= "000000";
                when "01101010011100" => rgb <= "000000";
                when "01101010011101" => rgb <= "000000";
                when "01101010011110" => rgb <= "000000";
                when "01101010011111" => rgb <= "000011";
                when "01101010100000" => rgb <= "000011";
                when "01101010100001" => rgb <= "000011";
                when "01101010100010" => rgb <= "000011";
                when "01101100000000" => rgb <= "000000";
                when "01101100000001" => rgb <= "000000";
                when "01101100000010" => rgb <= "000000";
                when "01101100000011" => rgb <= "000000";
                when "01101100000100" => rgb <= "000000";
                when "01101100000101" => rgb <= "000000";
                when "01101100000110" => rgb <= "000000";
                when "01101100000111" => rgb <= "000000";
                when "01101100001000" => rgb <= "000000";
                when "01101100001001" => rgb <= "000000";
                when "01101100001010" => rgb <= "000000";
                when "01101100001011" => rgb <= "000000";
                when "01101100001100" => rgb <= "000000";
                when "01101100001101" => rgb <= "000000";
                when "01101100001110" => rgb <= "000000";
                when "01101100001111" => rgb <= "000000";
                when "01101100010000" => rgb <= "000000";
                when "01101100010001" => rgb <= "000000";
                when "01101100010010" => rgb <= "000000";
                when "01101100010011" => rgb <= "000000";
                when "01101100010100" => rgb <= "000000";
                when "01101100010101" => rgb <= "000000";
                when "01101100010110" => rgb <= "000000";
                when "01101100010111" => rgb <= "000000";
                when "01101100011000" => rgb <= "000000";
                when "01101100011001" => rgb <= "000000";
                when "01101100011010" => rgb <= "000000";
                when "01101100011011" => rgb <= "000000";
                when "01101100011100" => rgb <= "000000";
                when "01101100011101" => rgb <= "000000";
                when "01101100011110" => rgb <= "000000";
                when "01101100011111" => rgb <= "000011";
                when "01101100100000" => rgb <= "000011";
                when "01101100100001" => rgb <= "000011";
                when "01101100100010" => rgb <= "000011";
                when "01101110000000" => rgb <= "000000";
                when "01101110000001" => rgb <= "000000";
                when "01101110000010" => rgb <= "000000";
                when "01101110000011" => rgb <= "000000";
                when "01101110000100" => rgb <= "000000";
                when "01101110000101" => rgb <= "000000";
                when "01101110000110" => rgb <= "000000";
                when "01101110000111" => rgb <= "000000";
                when "01101110001000" => rgb <= "000000";
                when "01101110001001" => rgb <= "000000";
                when "01101110001010" => rgb <= "000000";
                when "01101110001011" => rgb <= "000000";
                when "01101110001100" => rgb <= "000000";
                when "01101110001101" => rgb <= "000000";
                when "01101110001110" => rgb <= "000000";
                when "01101110001111" => rgb <= "000000";
                when "01101110010000" => rgb <= "000000";
                when "01101110010001" => rgb <= "000000";
                when "01101110010010" => rgb <= "000000";
                when "01101110010011" => rgb <= "000000";
                when "01101110010100" => rgb <= "000000";
                when "01101110010101" => rgb <= "000000";
                when "01101110010110" => rgb <= "000000";
                when "01101110010111" => rgb <= "000000";
                when "01101110011000" => rgb <= "000000";
                when "01101110011001" => rgb <= "000000";
                when "01101110011010" => rgb <= "000000";
                when "01101110011011" => rgb <= "000000";
                when "01101110011100" => rgb <= "000000";
                when "01101110011101" => rgb <= "000000";
                when "01101110011110" => rgb <= "000000";
                when "01101110011111" => rgb <= "000011";
                when "01101110100000" => rgb <= "000011";
                when "01101110100001" => rgb <= "000011";
                when "01101110100010" => rgb <= "000011";
                when "01110000000000" => rgb <= "000000";
                when "01110000000001" => rgb <= "000000";
                when "01110000000010" => rgb <= "000000";
                when "01110000000011" => rgb <= "000000";
                when "01110000000100" => rgb <= "000000";
                when "01110000000101" => rgb <= "000000";
                when "01110000000110" => rgb <= "000000";
                when "01110000000111" => rgb <= "000000";
                when "01110000001000" => rgb <= "000000";
                when "01110000001001" => rgb <= "000000";
                when "01110000001010" => rgb <= "000000";
                when "01110000001011" => rgb <= "000000";
                when "01110000001100" => rgb <= "000000";
                when "01110000001101" => rgb <= "000000";
                when "01110000001110" => rgb <= "000000";
                when "01110000001111" => rgb <= "000000";
                when "01110000010000" => rgb <= "000000";
                when "01110000010001" => rgb <= "000000";
                when "01110000010010" => rgb <= "000000";
                when "01110000010011" => rgb <= "000000";
                when "01110000010100" => rgb <= "000000";
                when "01110000010101" => rgb <= "000000";
                when "01110000010110" => rgb <= "000000";
                when "01110000010111" => rgb <= "000000";
                when "01110000011000" => rgb <= "000000";
                when "01110000011001" => rgb <= "000000";
                when "01110000011010" => rgb <= "000000";
                when "01110000011011" => rgb <= "000000";
                when "01110000011100" => rgb <= "000000";
                when "01110000011101" => rgb <= "000000";
                when "01110000011110" => rgb <= "000000";
                when "01110000011111" => rgb <= "000011";
                when "01110000100000" => rgb <= "000011";
                when "01110000100001" => rgb <= "000011";
                when "01110000100010" => rgb <= "000011";
                when "01110010000000" => rgb <= "000000";
                when "01110010000001" => rgb <= "000000";
                when "01110010000010" => rgb <= "000000";
                when "01110010000011" => rgb <= "000000";
                when "01110010000100" => rgb <= "000000";
                when "01110010000101" => rgb <= "000000";
                when "01110010000110" => rgb <= "000000";
                when "01110010000111" => rgb <= "000000";
                when "01110010001000" => rgb <= "000000";
                when "01110010001001" => rgb <= "000000";
                when "01110010001010" => rgb <= "000000";
                when "01110010001011" => rgb <= "000000";
                when "01110010001100" => rgb <= "000000";
                when "01110010001101" => rgb <= "000000";
                when "01110010001110" => rgb <= "000000";
                when "01110010001111" => rgb <= "000000";
                when "01110010010000" => rgb <= "000000";
                when "01110010010001" => rgb <= "000000";
                when "01110010010010" => rgb <= "000000";
                when "01110010010011" => rgb <= "000000";
                when "01110010010100" => rgb <= "000000";
                when "01110010010101" => rgb <= "000000";
                when "01110010010110" => rgb <= "000000";
                when "01110010010111" => rgb <= "000000";
                when "01110010011000" => rgb <= "000000";
                when "01110010011001" => rgb <= "000000";
                when "01110010011010" => rgb <= "000000";
                when "01110010011011" => rgb <= "000000";
                when "01110010011100" => rgb <= "000000";
                when "01110010011101" => rgb <= "000000";
                when "01110010011110" => rgb <= "000000";
                when "01110010011111" => rgb <= "000011";
                when "01110010100000" => rgb <= "000011";
                when "01110010100001" => rgb <= "000011";
                when "01110010100010" => rgb <= "000011";
                when "01110100000000" => rgb <= "000000";
                when "01110100000001" => rgb <= "000000";
                when "01110100000010" => rgb <= "000000";
                when "01110100000011" => rgb <= "000000";
                when "01110100000100" => rgb <= "000000";
                when "01110100000101" => rgb <= "000000";
                when "01110100000110" => rgb <= "000000";
                when "01110100000111" => rgb <= "000000";
                when "01110100001000" => rgb <= "000000";
                when "01110100001001" => rgb <= "000000";
                when "01110100001010" => rgb <= "000000";
                when "01110100001011" => rgb <= "000000";
                when "01110100001100" => rgb <= "000000";
                when "01110100001101" => rgb <= "000000";
                when "01110100001110" => rgb <= "000000";
                when "01110100001111" => rgb <= "000000";
                when "01110100010000" => rgb <= "000000";
                when "01110100010001" => rgb <= "000000";
                when "01110100010010" => rgb <= "000000";
                when "01110100010011" => rgb <= "000000";
                when "01110100010100" => rgb <= "000000";
                when "01110100010101" => rgb <= "000000";
                when "01110100010110" => rgb <= "000000";
                when "01110100010111" => rgb <= "000000";
                when "01110100011000" => rgb <= "000000";
                when "01110100011001" => rgb <= "000000";
                when "01110100011010" => rgb <= "000000";
                when "01110100011011" => rgb <= "000000";
                when "01110100011100" => rgb <= "000000";
                when "01110100011101" => rgb <= "000000";
                when "01110100011110" => rgb <= "000000";
                when "01110100011111" => rgb <= "000011";
                when "01110100100000" => rgb <= "000011";
                when "01110100100001" => rgb <= "000011";
                when "01110100100010" => rgb <= "000011";
                when "01110110000000" => rgb <= "000000";
                when "01110110000001" => rgb <= "000000";
                when "01110110000010" => rgb <= "000000";
                when "01110110000011" => rgb <= "000000";
                when "01110110000100" => rgb <= "000000";
                when "01110110000101" => rgb <= "000000";
                when "01110110000110" => rgb <= "000000";
                when "01110110000111" => rgb <= "000000";
                when "01110110001000" => rgb <= "000000";
                when "01110110001001" => rgb <= "000000";
                when "01110110001010" => rgb <= "000000";
                when "01110110001011" => rgb <= "000000";
                when "01110110001100" => rgb <= "000000";
                when "01110110001101" => rgb <= "000000";
                when "01110110001110" => rgb <= "000000";
                when "01110110001111" => rgb <= "000000";
                when "01110110010000" => rgb <= "000000";
                when "01110110010001" => rgb <= "000000";
                when "01110110010010" => rgb <= "000000";
                when "01110110010011" => rgb <= "000000";
                when "01110110010100" => rgb <= "000000";
                when "01110110010101" => rgb <= "000000";
                when "01110110010110" => rgb <= "000000";
                when "01110110010111" => rgb <= "000000";
                when "01110110011000" => rgb <= "000000";
                when "01110110011001" => rgb <= "000000";
                when "01110110011010" => rgb <= "000000";
                when "01110110011011" => rgb <= "000000";
                when "01110110011100" => rgb <= "000000";
                when "01110110011101" => rgb <= "000000";
                when "01110110011110" => rgb <= "000000";
                when "01110110011111" => rgb <= "000011";
                when "01110110100000" => rgb <= "000011";
                when "01110110100001" => rgb <= "000011";
                when "01110110100010" => rgb <= "000011";
                when "01111000000000" => rgb <= "000000";
                when "01111000000001" => rgb <= "000000";
                when "01111000000010" => rgb <= "000000";
                when "01111000000011" => rgb <= "000000";
                when "01111000000100" => rgb <= "000000";
                when "01111000000101" => rgb <= "000000";
                when "01111000000110" => rgb <= "000000";
                when "01111000000111" => rgb <= "000000";
                when "01111000001000" => rgb <= "000000";
                when "01111000001001" => rgb <= "000000";
                when "01111000001010" => rgb <= "000000";
                when "01111000001011" => rgb <= "000000";
                when "01111000001100" => rgb <= "000000";
                when "01111000001101" => rgb <= "000000";
                when "01111000001110" => rgb <= "000000";
                when "01111000001111" => rgb <= "000000";
                when "01111000010000" => rgb <= "000000";
                when "01111000010001" => rgb <= "000000";
                when "01111000010010" => rgb <= "000000";
                when "01111000010011" => rgb <= "000000";
                when "01111000010100" => rgb <= "000000";
                when "01111000010101" => rgb <= "000000";
                when "01111000010110" => rgb <= "000000";
                when "01111000010111" => rgb <= "000000";
                when "01111000011000" => rgb <= "000000";
                when "01111000011001" => rgb <= "000000";
                when "01111000011010" => rgb <= "000000";
                when "01111000011011" => rgb <= "000000";
                when "01111000011100" => rgb <= "000000";
                when "01111000011101" => rgb <= "000000";
                when "01111000011110" => rgb <= "000000";
                when "01111000011111" => rgb <= "000011";
                when "01111000100000" => rgb <= "000011";
                when "01111000100001" => rgb <= "000011";
                when "01111000100010" => rgb <= "000011";
                when "01111010000000" => rgb <= "000000";
                when "01111010000001" => rgb <= "000000";
                when "01111010000010" => rgb <= "000000";
                when "01111010000011" => rgb <= "000000";
                when "01111010000100" => rgb <= "000000";
                when "01111010000101" => rgb <= "000000";
                when "01111010000110" => rgb <= "000000";
                when "01111010000111" => rgb <= "000000";
                when "01111010001000" => rgb <= "000000";
                when "01111010001001" => rgb <= "000000";
                when "01111010001010" => rgb <= "000000";
                when "01111010001011" => rgb <= "000000";
                when "01111010001100" => rgb <= "000000";
                when "01111010001101" => rgb <= "000000";
                when "01111010001110" => rgb <= "000000";
                when "01111010001111" => rgb <= "000000";
                when "01111010010000" => rgb <= "000000";
                when "01111010010001" => rgb <= "000000";
                when "01111010010010" => rgb <= "000000";
                when "01111010010011" => rgb <= "000000";
                when "01111010010100" => rgb <= "000000";
                when "01111010010101" => rgb <= "000000";
                when "01111010010110" => rgb <= "000000";
                when "01111010010111" => rgb <= "000000";
                when "01111010011000" => rgb <= "000000";
                when "01111010011001" => rgb <= "000000";
                when "01111010011010" => rgb <= "000000";
                when "01111010011011" => rgb <= "000000";
                when "01111010011100" => rgb <= "000000";
                when "01111010011101" => rgb <= "000000";
                when "01111010011110" => rgb <= "000000";
                when "01111010011111" => rgb <= "000011";
                when "01111010100000" => rgb <= "000011";
                when "01111010100001" => rgb <= "000011";
                when "01111010100010" => rgb <= "000011";
                when "01111100000000" => rgb <= "000000";
                when "01111100000001" => rgb <= "000000";
                when "01111100000010" => rgb <= "000000";
                when "01111100000011" => rgb <= "000000";
                when "01111100000100" => rgb <= "000000";
                when "01111100000101" => rgb <= "000000";
                when "01111100000110" => rgb <= "000000";
                when "01111100000111" => rgb <= "000000";
                when "01111100001000" => rgb <= "000000";
                when "01111100001001" => rgb <= "000000";
                when "01111100001010" => rgb <= "000000";
                when "01111100001011" => rgb <= "000000";
                when "01111100001100" => rgb <= "000000";
                when "01111100001101" => rgb <= "000000";
                when "01111100001110" => rgb <= "000000";
                when "01111100001111" => rgb <= "000000";
                when "01111100010000" => rgb <= "000000";
                when "01111100010001" => rgb <= "000000";
                when "01111100010010" => rgb <= "000000";
                when "01111100010011" => rgb <= "000000";
                when "01111100010100" => rgb <= "000000";
                when "01111100010101" => rgb <= "000000";
                when "01111100010110" => rgb <= "000000";
                when "01111100010111" => rgb <= "000000";
                when "01111100011000" => rgb <= "000000";
                when "01111100011001" => rgb <= "000000";
                when "01111100011010" => rgb <= "000000";
                when "01111100011011" => rgb <= "000000";
                when "01111100011100" => rgb <= "000000";
                when "01111100011101" => rgb <= "000000";
                when "01111100011110" => rgb <= "000000";
                when "01111100011111" => rgb <= "000011";
                when "01111100100000" => rgb <= "000011";
                when "01111100100001" => rgb <= "000011";
                when "01111100100010" => rgb <= "000011";
                when "01111110000000" => rgb <= "000000";
                when "01111110000001" => rgb <= "000000";
                when "01111110000010" => rgb <= "000000";
                when "01111110000011" => rgb <= "000000";
                when "01111110000100" => rgb <= "000000";
                when "01111110000101" => rgb <= "000000";
                when "01111110000110" => rgb <= "000000";
                when "01111110000111" => rgb <= "000000";
                when "01111110001000" => rgb <= "000000";
                when "01111110001001" => rgb <= "000000";
                when "01111110001010" => rgb <= "000000";
                when "01111110001011" => rgb <= "000000";
                when "01111110001100" => rgb <= "000000";
                when "01111110001101" => rgb <= "000000";
                when "01111110001110" => rgb <= "000000";
                when "01111110001111" => rgb <= "000000";
                when "01111110010000" => rgb <= "000000";
                when "01111110010001" => rgb <= "000000";
                when "01111110010010" => rgb <= "000000";
                when "01111110010011" => rgb <= "000000";
                when "01111110010100" => rgb <= "000000";
                when "01111110010101" => rgb <= "000000";
                when "01111110010110" => rgb <= "000000";
                when "01111110010111" => rgb <= "000000";
                when "01111110011000" => rgb <= "000000";
                when "01111110011001" => rgb <= "000000";
                when "01111110011010" => rgb <= "000000";
                when "01111110011011" => rgb <= "000000";
                when "01111110011100" => rgb <= "000000";
                when "01111110011101" => rgb <= "000000";
                when "01111110011110" => rgb <= "000000";
                when "01111110011111" => rgb <= "000011";
                when "01111110100000" => rgb <= "000011";
                when "01111110100001" => rgb <= "000011";
                when "01111110100010" => rgb <= "000011";
                when "10000000000000" => rgb <= "000000";
                when "10000000000001" => rgb <= "000000";
                when "10000000000010" => rgb <= "000000";
                when "10000000000011" => rgb <= "000000";
                when "10000000000100" => rgb <= "000000";
                when "10000000000101" => rgb <= "000000";
                when "10000000000110" => rgb <= "000000";
                when "10000000000111" => rgb <= "000000";
                when "10000000001000" => rgb <= "000000";
                when "10000000001001" => rgb <= "000000";
                when "10000000001010" => rgb <= "000000";
                when "10000000001011" => rgb <= "000000";
                when "10000000001100" => rgb <= "000000";
                when "10000000001101" => rgb <= "000000";
                when "10000000001110" => rgb <= "000000";
                when "10000000001111" => rgb <= "000000";
                when "10000000010000" => rgb <= "000000";
                when "10000000010001" => rgb <= "000000";
                when "10000000010010" => rgb <= "000000";
                when "10000000010011" => rgb <= "000000";
                when "10000000010100" => rgb <= "000000";
                when "10000000010101" => rgb <= "000000";
                when "10000000010110" => rgb <= "000000";
                when "10000000010111" => rgb <= "000000";
                when "10000000011000" => rgb <= "000000";
                when "10000000011001" => rgb <= "000000";
                when "10000000011010" => rgb <= "000000";
                when "10000000011011" => rgb <= "000000";
                when "10000000011100" => rgb <= "000000";
                when "10000000011101" => rgb <= "000000";
                when "10000000011110" => rgb <= "000000";
                when "10000000011111" => rgb <= "000011";
                when "10000000100000" => rgb <= "000011";
                when "10000000100001" => rgb <= "000011";
                when "10000000100010" => rgb <= "000011";
                when "10000010000000" => rgb <= "000000";
                when "10000010000001" => rgb <= "000000";
                when "10000010000010" => rgb <= "000000";
                when "10000010000011" => rgb <= "000000";
                when "10000010000100" => rgb <= "000000";
                when "10000010000101" => rgb <= "000000";
                when "10000010000110" => rgb <= "000000";
                when "10000010000111" => rgb <= "000000";
                when "10000010001000" => rgb <= "000000";
                when "10000010001001" => rgb <= "000000";
                when "10000010001010" => rgb <= "000000";
                when "10000010001011" => rgb <= "000000";
                when "10000010001100" => rgb <= "000000";
                when "10000010001101" => rgb <= "000000";
                when "10000010001110" => rgb <= "000000";
                when "10000010001111" => rgb <= "000000";
                when "10000010010000" => rgb <= "000000";
                when "10000010010001" => rgb <= "000000";
                when "10000010010010" => rgb <= "000000";
                when "10000010010011" => rgb <= "000000";
                when "10000010010100" => rgb <= "000000";
                when "10000010010101" => rgb <= "000000";
                when "10000010010110" => rgb <= "000000";
                when "10000010010111" => rgb <= "000000";
                when "10000010011000" => rgb <= "000000";
                when "10000010011001" => rgb <= "000000";
                when "10000010011010" => rgb <= "000000";
                when "10000010011011" => rgb <= "000000";
                when "10000010011100" => rgb <= "000000";
                when "10000010011101" => rgb <= "000000";
                when "10000010011110" => rgb <= "000000";
                when "10000010011111" => rgb <= "000011";
                when "10000010100000" => rgb <= "000011";
                when "10000010100001" => rgb <= "000011";
                when "10000010100010" => rgb <= "000011";
                when "10000100000000" => rgb <= "000000";
                when "10000100000001" => rgb <= "000000";
                when "10000100000010" => rgb <= "000000";
                when "10000100000011" => rgb <= "000000";
                when "10000100000100" => rgb <= "000000";
                when "10000100000101" => rgb <= "000000";
                when "10000100000110" => rgb <= "000000";
                when "10000100000111" => rgb <= "000000";
                when "10000100001000" => rgb <= "000000";
                when "10000100001001" => rgb <= "000000";
                when "10000100001010" => rgb <= "000000";
                when "10000100001011" => rgb <= "000000";
                when "10000100001100" => rgb <= "000000";
                when "10000100001101" => rgb <= "000000";
                when "10000100001110" => rgb <= "000000";
                when "10000100001111" => rgb <= "000000";
                when "10000100010000" => rgb <= "000000";
                when "10000100010001" => rgb <= "000000";
                when "10000100010010" => rgb <= "000000";
                when "10000100010011" => rgb <= "000000";
                when "10000100010100" => rgb <= "000000";
                when "10000100010101" => rgb <= "000000";
                when "10000100010110" => rgb <= "000000";
                when "10000100010111" => rgb <= "000000";
                when "10000100011000" => rgb <= "000000";
                when "10000100011001" => rgb <= "000000";
                when "10000100011010" => rgb <= "000000";
                when "10000100011011" => rgb <= "000000";
                when "10000100011100" => rgb <= "000000";
                when "10000100011101" => rgb <= "000000";
                when "10000100011110" => rgb <= "000000";
                when "10000100011111" => rgb <= "000011";
                when "10000100100000" => rgb <= "000011";
                when "10000100100001" => rgb <= "000011";
                when "10000100100010" => rgb <= "000011";
                when "10000110000000" => rgb <= "000000";
                when "10000110000001" => rgb <= "000000";
                when "10000110000010" => rgb <= "000000";
                when "10000110000011" => rgb <= "000000";
                when "10000110000100" => rgb <= "000000";
                when "10000110000101" => rgb <= "000000";
                when "10000110000110" => rgb <= "000000";
                when "10000110000111" => rgb <= "000000";
                when "10000110001000" => rgb <= "000000";
                when "10000110001001" => rgb <= "000000";
                when "10000110001010" => rgb <= "000000";
                when "10000110001011" => rgb <= "000000";
                when "10000110001100" => rgb <= "000000";
                when "10000110001101" => rgb <= "000000";
                when "10000110001110" => rgb <= "000000";
                when "10000110001111" => rgb <= "000000";
                when "10000110010000" => rgb <= "000000";
                when "10000110010001" => rgb <= "000000";
                when "10000110010010" => rgb <= "000000";
                when "10000110010011" => rgb <= "000000";
                when "10000110010100" => rgb <= "000000";
                when "10000110010101" => rgb <= "000000";
                when "10000110010110" => rgb <= "000000";
                when "10000110010111" => rgb <= "000000";
                when "10000110011000" => rgb <= "000000";
                when "10000110011001" => rgb <= "000000";
                when "10000110011010" => rgb <= "000000";
                when "10000110011011" => rgb <= "000000";
                when "10000110011100" => rgb <= "000000";
                when "10000110011101" => rgb <= "000000";
                when "10000110011110" => rgb <= "000000";
                when "10000110011111" => rgb <= "000011";
                when "10000110100000" => rgb <= "000011";
                when "10000110100001" => rgb <= "000011";
                when "10000110100010" => rgb <= "000011";
                when "10001000000000" => rgb <= "000000";
                when "10001000000001" => rgb <= "000000";
                when "10001000000010" => rgb <= "000000";
                when "10001000000011" => rgb <= "000000";
                when "10001000000100" => rgb <= "000000";
                when "10001000000101" => rgb <= "000000";
                when "10001000000110" => rgb <= "000000";
                when "10001000000111" => rgb <= "000000";
                when "10001000001000" => rgb <= "000000";
                when "10001000001001" => rgb <= "000000";
                when "10001000001010" => rgb <= "000000";
                when "10001000001011" => rgb <= "000000";
                when "10001000001100" => rgb <= "000000";
                when "10001000001101" => rgb <= "000000";
                when "10001000001110" => rgb <= "000000";
                when "10001000001111" => rgb <= "000000";
                when "10001000010000" => rgb <= "000000";
                when "10001000010001" => rgb <= "000000";
                when "10001000010010" => rgb <= "000000";
                when "10001000010011" => rgb <= "000000";
                when "10001000010100" => rgb <= "000000";
                when "10001000010101" => rgb <= "000000";
                when "10001000010110" => rgb <= "000000";
                when "10001000010111" => rgb <= "000000";
                when "10001000011000" => rgb <= "000000";
                when "10001000011001" => rgb <= "000000";
                when "10001000011010" => rgb <= "000000";
                when "10001000011011" => rgb <= "000000";
                when "10001000011100" => rgb <= "000000";
                when "10001000011101" => rgb <= "000000";
                when "10001000011110" => rgb <= "000000";
                when "10001000011111" => rgb <= "000011";
                when "10001000100000" => rgb <= "000011";
                when "10001000100001" => rgb <= "000011";
                when "10001000100010" => rgb <= "000011";
                when "10001010000000" => rgb <= "000000";
                when "10001010000001" => rgb <= "000000";
                when "10001010000010" => rgb <= "000000";
                when "10001010000011" => rgb <= "000000";
                when "10001010000100" => rgb <= "000000";
                when "10001010000101" => rgb <= "000000";
                when "10001010000110" => rgb <= "000000";
                when "10001010000111" => rgb <= "000000";
                when "10001010001000" => rgb <= "000000";
                when "10001010001001" => rgb <= "000000";
                when "10001010001010" => rgb <= "000000";
                when "10001010001011" => rgb <= "000000";
                when "10001010001100" => rgb <= "000000";
                when "10001010001101" => rgb <= "000000";
                when "10001010001110" => rgb <= "000000";
                when "10001010001111" => rgb <= "000000";
                when "10001010010000" => rgb <= "000000";
                when "10001010010001" => rgb <= "000000";
                when "10001010010010" => rgb <= "000000";
                when "10001010010011" => rgb <= "000000";
                when "10001010010100" => rgb <= "000000";
                when "10001010010101" => rgb <= "000000";
                when "10001010010110" => rgb <= "000000";
                when "10001010010111" => rgb <= "000000";
                when "10001010011000" => rgb <= "000000";
                when "10001010011001" => rgb <= "000000";
                when "10001010011010" => rgb <= "000000";
                when "10001010011011" => rgb <= "000000";
                when "10001010011100" => rgb <= "000000";
                when "10001010011101" => rgb <= "000000";
                when "10001010011110" => rgb <= "000000";
                when "10001010011111" => rgb <= "000011";
                when "10001010100000" => rgb <= "000011";
                when "10001010100001" => rgb <= "000011";
                when "10001010100010" => rgb <= "000011";
                when others => rgb <= "111111";
               
                end case;
            end if;
            end process;
        end;
                
