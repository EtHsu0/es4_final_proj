library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gapple is
    port (
        row : in unsigned (9 downto 0);
        col : in unsigned (9 downto 0);
        clk : in std_logic;
        rgb : out unsigned(5 downto 0)
    );
end gapple;

architecture synth of gapple is
    signal addr : unsigned(11 downto 0);

    begin
        addr <= unsigned(row(5 downto 0)) & unsigned(col(5 downto 0));
        process(clk) is begin
            if rising_edge(clk) then
				if (row(9 downto 6) = "00000" and col(9 downto 6) = "00000") then			
                case addr is 
                          when "000000000000" => rgb <= "000000";
                          when "000000000001" => rgb <= "000000";
                          when "000000000010" => rgb <= "000000";
                          when "000000000011" => rgb <= "000000";
                          when "000000000100" => rgb <= "000000";
                          when "000000000101" => rgb <= "000000";
                          when "000000000110" => rgb <= "000000";
                          when "000000000111" => rgb <= "000000";
                          when "000000001000" => rgb <= "000000";
                          when "000000001001" => rgb <= "000000";
                          when "000000001010" => rgb <= "000000";
                          when "000000001011" => rgb <= "000000";
                          when "000000001100" => rgb <= "000000";
                          when "000000001101" => rgb <= "000000";
                          when "000000001110" => rgb <= "000000";
                          when "000000001111" => rgb <= "000000";
                          when "000000010000" => rgb <= "000000";
                          when "000000010001" => rgb <= "000000";
                          when "000000010010" => rgb <= "000000";
                          when "000000010011" => rgb <= "000000";
                          when "000000010100" => rgb <= "000000";
                          when "000000010101" => rgb <= "000000";
                          when "000000010110" => rgb <= "000000";
                          when "000000010111" => rgb <= "000000";
                          when "000000011000" => rgb <= "000000";
                          when "000000011001" => rgb <= "000000";
                          when "000000011010" => rgb <= "000000";
                          when "000000011011" => rgb <= "000000";
                          when "000000011100" => rgb <= "000000";
                          when "000000011101" => rgb <= "000000";
                          when "000000011110" => rgb <= "000000";
                          when "000000011111" => rgb <= "000000";
                          when "000000100000" => rgb <= "000000";
                          when "000000100001" => rgb <= "000000";
                          when "000000100010" => rgb <= "000000";
                          when "000000100011" => rgb <= "000000";
                          when "000000100100" => rgb <= "000000";
                          when "000000100101" => rgb <= "000000";
                          when "000000100110" => rgb <= "000000";
                          when "000000100111" => rgb <= "000000";
                          when "000000101000" => rgb <= "000000";
                          when "000000101001" => rgb <= "000000";
                          when "000001000000" => rgb <= "000000";
                          when "000001000001" => rgb <= "000000";
                          when "000001000010" => rgb <= "000000";
                          when "000001000011" => rgb <= "000000";
                          when "000001000100" => rgb <= "000000";
                          when "000001000101" => rgb <= "000000";
                          when "000001000110" => rgb <= "000000";
                          when "000001000111" => rgb <= "000000";
                          when "000001001000" => rgb <= "000000";
                          when "000001001001" => rgb <= "000000";
                          when "000001001010" => rgb <= "000000";
                          when "000001001011" => rgb <= "000000";
                          when "000001001100" => rgb <= "000000";
                          when "000001001101" => rgb <= "000000";
                          when "000001001110" => rgb <= "000000";
                          when "000001001111" => rgb <= "000000";
                          when "000001010000" => rgb <= "000000";
                          when "000001010001" => rgb <= "000000";
                          when "000001010010" => rgb <= "000000";
                          when "000001010011" => rgb <= "000000";
                          when "000001010100" => rgb <= "000000";
                          when "000001010101" => rgb <= "000000";
                          when "000001010110" => rgb <= "000000";
                          when "000001010111" => rgb <= "000000";
                          when "000001011000" => rgb <= "001000";
                          when "000001011001" => rgb <= "001000";
                          when "000001011010" => rgb <= "001000";
                          when "000001011011" => rgb <= "001000";
                          when "000001011100" => rgb <= "001000";
                          when "000001011101" => rgb <= "001000";
                          when "000001011110" => rgb <= "001000";
                          when "000001011111" => rgb <= "001000";
                          when "000001100000" => rgb <= "000000";
                          when "000001100001" => rgb <= "000000";
                          when "000001100010" => rgb <= "000000";
                          when "000001100011" => rgb <= "000000";
                          when "000001100100" => rgb <= "000000";
                          when "000001100101" => rgb <= "000000";
                          when "000001100110" => rgb <= "000000";
                          when "000001100111" => rgb <= "000000";
                          when "000001101000" => rgb <= "000000";
                          when "000001101001" => rgb <= "000000";
                          when "000010000000" => rgb <= "000000";
                          when "000010000001" => rgb <= "000000";
                          when "000010000010" => rgb <= "000000";
                          when "000010000011" => rgb <= "000000";
                          when "000010000100" => rgb <= "000000";
                          when "000010000101" => rgb <= "000000";
                          when "000010000110" => rgb <= "000000";
                          when "000010000111" => rgb <= "000000";
                          when "000010001000" => rgb <= "000000";
                          when "000010001001" => rgb <= "000000";
                          when "000010001010" => rgb <= "000000";
                          when "000010001011" => rgb <= "000000";
                          when "000010001100" => rgb <= "000000";
                          when "000010001101" => rgb <= "000000";
                          when "000010001110" => rgb <= "000000";
                          when "000010001111" => rgb <= "000000";
                          when "000010010000" => rgb <= "000000";
                          when "000010010001" => rgb <= "000000";
                          when "000010010010" => rgb <= "000000";
                          when "000010010011" => rgb <= "000000";
                          when "000010010100" => rgb <= "000000";
                          when "000010010101" => rgb <= "000000";
                          when "000010010110" => rgb <= "000000";
                          when "000010010111" => rgb <= "000000";
                          when "000010011000" => rgb <= "001000";
                          when "000010011001" => rgb <= "001000";
                          when "000010011010" => rgb <= "001000";
                          when "000010011011" => rgb <= "001000";
                          when "000010011100" => rgb <= "001000";
                          when "000010011101" => rgb <= "001000";
                          when "000010011110" => rgb <= "001000";
                          when "000010011111" => rgb <= "001000";
                          when "000010100000" => rgb <= "000000";
                          when "000010100001" => rgb <= "000000";
                          when "000010100010" => rgb <= "000000";
                          when "000010100011" => rgb <= "000000";
                          when "000010100100" => rgb <= "000000";
                          when "000010100101" => rgb <= "000000";
                          when "000010100110" => rgb <= "000000";
                          when "000010100111" => rgb <= "000000";
                          when "000010101000" => rgb <= "000000";
                          when "000010101001" => rgb <= "000000";
                          when "000011000000" => rgb <= "000000";
                          when "000011000001" => rgb <= "000000";
                          when "000011000010" => rgb <= "000000";
                          when "000011000011" => rgb <= "000000";
                          when "000011000100" => rgb <= "000000";
                          when "000011000101" => rgb <= "000000";
                          when "000011000110" => rgb <= "000000";
                          when "000011000111" => rgb <= "000000";
                          when "000011001000" => rgb <= "000000";
                          when "000011001001" => rgb <= "000000";
                          when "000011001010" => rgb <= "000000";
                          when "000011001011" => rgb <= "000000";
                          when "000011001100" => rgb <= "000000";
                          when "000011001101" => rgb <= "000000";
                          when "000011001110" => rgb <= "000000";
                          when "000011001111" => rgb <= "000000";
                          when "000011010000" => rgb <= "000000";
                          when "000011010001" => rgb <= "000000";
                          when "000011010010" => rgb <= "000000";
                          when "000011010011" => rgb <= "000000";
                          when "000011010100" => rgb <= "000000";
                          when "000011010101" => rgb <= "000000";
                          when "000011010110" => rgb <= "000000";
                          when "000011010111" => rgb <= "001000";
                          when "000011011000" => rgb <= "001000";
                          when "000011011001" => rgb <= "001000";
                          when "000011011010" => rgb <= "001000";
                          when "000011011011" => rgb <= "001000";
                          when "000011011100" => rgb <= "001000";
                          when "000011011101" => rgb <= "001000";
                          when "000011011110" => rgb <= "001000";
                          when "000011011111" => rgb <= "001000";
                          when "000011100000" => rgb <= "001000";
                          when "000011100001" => rgb <= "001000";
                          when "000011100010" => rgb <= "000000";
                          when "000011100011" => rgb <= "000000";
                          when "000011100100" => rgb <= "000000";
                          when "000011100101" => rgb <= "000000";
                          when "000011100110" => rgb <= "000000";
                          when "000011100111" => rgb <= "000000";
                          when "000011101000" => rgb <= "000000";
                          when "000011101001" => rgb <= "000000";
                          when "000100000000" => rgb <= "000000";
                          when "000100000001" => rgb <= "000000";
                          when "000100000010" => rgb <= "000000";
                          when "000100000011" => rgb <= "000000";
                          when "000100000100" => rgb <= "000000";
                          when "000100000101" => rgb <= "000000";
                          when "000100000110" => rgb <= "000000";
                          when "000100000111" => rgb <= "000000";
                          when "000100001000" => rgb <= "000000";
                          when "000100001001" => rgb <= "000000";
                          when "000100001010" => rgb <= "000000";
                          when "000100001011" => rgb <= "000000";
                          when "000100001100" => rgb <= "000000";
                          when "000100001101" => rgb <= "000000";
                          when "000100001110" => rgb <= "000000";
                          when "000100001111" => rgb <= "000000";
                          when "000100010000" => rgb <= "000000";
                          when "000100010001" => rgb <= "000000";
                          when "000100010010" => rgb <= "000000";
                          when "000100010011" => rgb <= "000000";
                          when "000100010100" => rgb <= "000000";
                          when "000100010101" => rgb <= "000000";
                          when "000100010110" => rgb <= "000000";
                          when "000100010111" => rgb <= "001000";
                          when "000100011000" => rgb <= "001000";
                          when "000100011001" => rgb <= "001000";
                          when "000100011010" => rgb <= "001000";
                          when "000100011011" => rgb <= "001000";
                          when "000100011100" => rgb <= "001000";
                          when "000100011101" => rgb <= "001000";
                          when "000100011110" => rgb <= "001000";
                          when "000100011111" => rgb <= "001000";
                          when "000100100000" => rgb <= "001000";
                          when "000100100001" => rgb <= "001000";
                          when "000100100010" => rgb <= "000000";
                          when "000100100011" => rgb <= "000000";
                          when "000100100100" => rgb <= "000000";
                          when "000100100101" => rgb <= "000000";
                          when "000100100110" => rgb <= "000000";
                          when "000100100111" => rgb <= "000000";
                          when "000100101000" => rgb <= "000000";
                          when "000100101001" => rgb <= "000000";
                          when "000101000000" => rgb <= "000000";
                          when "000101000001" => rgb <= "000000";
                          when "000101000010" => rgb <= "000000";
                          when "000101000011" => rgb <= "000000";
                          when "000101000100" => rgb <= "000000";
                          when "000101000101" => rgb <= "000000";
                          when "000101000110" => rgb <= "000000";
                          when "000101000111" => rgb <= "000000";
                          when "000101001000" => rgb <= "000000";
                          when "000101001001" => rgb <= "000000";
                          when "000101001010" => rgb <= "000000";
                          when "000101001011" => rgb <= "000000";
                          when "000101001100" => rgb <= "000000";
                          when "000101001101" => rgb <= "000000";
                          when "000101001110" => rgb <= "000000";
                          when "000101001111" => rgb <= "000000";
                          when "000101010000" => rgb <= "000000";
                          when "000101010001" => rgb <= "010000";
                          when "000101010010" => rgb <= "010000";
                          when "000101010011" => rgb <= "010000";
                          when "000101010100" => rgb <= "010000";
                          when "000101010101" => rgb <= "000000";
                          when "000101010110" => rgb <= "000000";
                          when "000101010111" => rgb <= "001000";
                          when "000101011000" => rgb <= "001000";
                          when "000101011001" => rgb <= "001000";
                          when "000101011010" => rgb <= "001000";
                          when "000101011011" => rgb <= "001000";
                          when "000101011100" => rgb <= "001000";
                          when "000101011101" => rgb <= "001000";
                          when "000101011110" => rgb <= "001000";
                          when "000101011111" => rgb <= "001000";
                          when "000101100000" => rgb <= "001000";
                          when "000101100001" => rgb <= "001000";
                          when "000101100010" => rgb <= "000000";
                          when "000101100011" => rgb <= "000000";
                          when "000101100100" => rgb <= "000000";
                          when "000101100101" => rgb <= "000000";
                          when "000101100110" => rgb <= "000000";
                          when "000101100111" => rgb <= "000000";
                          when "000101101000" => rgb <= "000000";
                          when "000101101001" => rgb <= "000000";
                          when "000110000000" => rgb <= "000000";
                          when "000110000001" => rgb <= "000000";
                          when "000110000010" => rgb <= "000000";
                          when "000110000011" => rgb <= "000000";
                          when "000110000100" => rgb <= "000000";
                          when "000110000101" => rgb <= "000000";
                          when "000110000110" => rgb <= "000000";
                          when "000110000111" => rgb <= "000000";
                          when "000110001000" => rgb <= "000000";
                          when "000110001001" => rgb <= "000000";
                          when "000110001010" => rgb <= "000000";
                          when "000110001011" => rgb <= "000000";
                          when "000110001100" => rgb <= "000000";
                          when "000110001101" => rgb <= "000000";
                          when "000110001110" => rgb <= "000000";
                          when "000110001111" => rgb <= "000000";
                          when "000110010000" => rgb <= "000000";
                          when "000110010001" => rgb <= "010000";
                          when "000110010010" => rgb <= "010000";
                          when "000110010011" => rgb <= "010000";
                          when "000110010100" => rgb <= "010000";
                          when "000110010101" => rgb <= "010000";
                          when "000110010110" => rgb <= "010000";
                          when "000110010111" => rgb <= "001000";
                          when "000110011000" => rgb <= "001000";
                          when "000110011001" => rgb <= "001000";
                          when "000110011010" => rgb <= "001000";
                          when "000110011011" => rgb <= "001000";
                          when "000110011100" => rgb <= "000000";
                          when "000110011101" => rgb <= "000000";
                          when "000110011110" => rgb <= "000000";
                          when "000110011111" => rgb <= "000000";
                          when "000110100000" => rgb <= "000000";
                          when "000110100001" => rgb <= "000000";
                          when "000110100010" => rgb <= "000000";
                          when "000110100011" => rgb <= "000000";
                          when "000110100100" => rgb <= "000000";
                          when "000110100101" => rgb <= "000000";
                          when "000110100110" => rgb <= "000000";
                          when "000110100111" => rgb <= "000000";
                          when "000110101000" => rgb <= "000000";
                          when "000110101001" => rgb <= "000000";
                          when "000111000000" => rgb <= "000000";
                          when "000111000001" => rgb <= "000000";
                          when "000111000010" => rgb <= "000000";
                          when "000111000011" => rgb <= "000000";
                          when "000111000100" => rgb <= "000000";
                          when "000111000101" => rgb <= "000000";
                          when "000111000110" => rgb <= "000000";
                          when "000111000111" => rgb <= "000000";
                          when "000111001000" => rgb <= "000000";
                          when "000111001001" => rgb <= "000000";
                          when "000111001010" => rgb <= "000000";
                          when "000111001011" => rgb <= "000000";
                          when "000111001100" => rgb <= "000000";
                          when "000111001101" => rgb <= "000000";
                          when "000111001110" => rgb <= "000000";
                          when "000111001111" => rgb <= "000000";
                          when "000111010000" => rgb <= "000000";
                          when "000111010001" => rgb <= "010000";
                          when "000111010010" => rgb <= "010000";
                          when "000111010011" => rgb <= "010000";
                          when "000111010100" => rgb <= "010000";
                          when "000111010101" => rgb <= "010000";
                          when "000111010110" => rgb <= "010000";
                          when "000111010111" => rgb <= "001000";
                          when "000111011000" => rgb <= "001000";
                          when "000111011001" => rgb <= "000000";
                          when "000111011010" => rgb <= "000000";
                          when "000111011011" => rgb <= "000000";
                          when "000111011100" => rgb <= "000000";
                          when "000111011101" => rgb <= "000000";
                          when "000111011110" => rgb <= "000000";
                          when "000111011111" => rgb <= "000000";
                          when "000111100000" => rgb <= "000000";
                          when "000111100001" => rgb <= "000000";
                          when "000111100010" => rgb <= "000000";
                          when "000111100011" => rgb <= "000000";
                          when "000111100100" => rgb <= "000000";
                          when "000111100101" => rgb <= "000000";
                          when "000111100110" => rgb <= "000000";
                          when "000111100111" => rgb <= "000000";
                          when "000111101000" => rgb <= "000000";
                          when "000111101001" => rgb <= "000000";
                          when "001000000000" => rgb <= "000000";
                          when "001000000001" => rgb <= "000000";
                          when "001000000010" => rgb <= "000000";
                          when "001000000011" => rgb <= "000000";
                          when "001000000100" => rgb <= "000000";
                          when "001000000101" => rgb <= "000000";
                          when "001000000110" => rgb <= "000000";
                          when "001000000111" => rgb <= "000000";
                          when "001000001000" => rgb <= "101000";
                          when "001000001001" => rgb <= "101000";
                          when "001000001010" => rgb <= "101000";
                          when "001000001011" => rgb <= "101000";
                          when "001000001100" => rgb <= "101000";
                          when "001000001101" => rgb <= "101000";
                          when "001000001110" => rgb <= "101000";
                          when "001000001111" => rgb <= "101000";
                          when "001000010000" => rgb <= "101000";
                          when "001000010001" => rgb <= "010100";
                          when "001000010010" => rgb <= "010000";
                          when "001000010011" => rgb <= "010000";
                          when "001000010100" => rgb <= "010000";
                          when "001000010101" => rgb <= "010000";
                          when "001000010110" => rgb <= "010000";
                          when "001000010111" => rgb <= "001000";
                          when "001000011000" => rgb <= "001000";
                          when "001000011001" => rgb <= "101000";
                          when "001000011010" => rgb <= "101000";
                          when "001000011011" => rgb <= "101000";
                          when "001000011100" => rgb <= "101000";
                          when "001000011101" => rgb <= "101000";
                          when "001000011110" => rgb <= "101000";
                          when "001000011111" => rgb <= "101000";
                          when "001000100000" => rgb <= "101000";
                          when "001000100001" => rgb <= "101000";
                          when "001000100010" => rgb <= "000000";
                          when "001000100011" => rgb <= "000000";
                          when "001000100100" => rgb <= "000000";
                          when "001000100101" => rgb <= "000000";
                          when "001000100110" => rgb <= "000000";
                          when "001000100111" => rgb <= "000000";
                          when "001000101000" => rgb <= "000000";
                          when "001000101001" => rgb <= "000000";
                          when "001001000000" => rgb <= "000000";
                          when "001001000001" => rgb <= "000000";
                          when "001001000010" => rgb <= "000000";
                          when "001001000011" => rgb <= "000000";
                          when "001001000100" => rgb <= "000000";
                          when "001001000101" => rgb <= "000000";
                          when "001001000110" => rgb <= "000000";
                          when "001001000111" => rgb <= "000000";
                          when "001001001000" => rgb <= "101000";
                          when "001001001001" => rgb <= "101000";
                          when "001001001010" => rgb <= "101000";
                          when "001001001011" => rgb <= "101000";
                          when "001001001100" => rgb <= "101000";
                          when "001001001101" => rgb <= "101000";
                          when "001001001110" => rgb <= "101000";
                          when "001001001111" => rgb <= "101000";
                          when "001001010000" => rgb <= "101000";
                          when "001001010001" => rgb <= "101000";
                          when "001001010010" => rgb <= "010000";
                          when "001001010011" => rgb <= "010000";
                          when "001001010100" => rgb <= "010000";
                          when "001001010101" => rgb <= "010000";
                          when "001001010110" => rgb <= "010000";
                          when "001001010111" => rgb <= "010000";
                          when "001001011000" => rgb <= "101000";
                          when "001001011001" => rgb <= "101000";
                          when "001001011010" => rgb <= "101000";
                          when "001001011011" => rgb <= "101000";
                          when "001001011100" => rgb <= "101000";
                          when "001001011101" => rgb <= "101000";
                          when "001001011110" => rgb <= "101000";
                          when "001001011111" => rgb <= "101000";
                          when "001001100000" => rgb <= "101000";
                          when "001001100001" => rgb <= "101000";
                          when "001001100010" => rgb <= "000000";
                          when "001001100011" => rgb <= "000000";
                          when "001001100100" => rgb <= "000000";
                          when "001001100101" => rgb <= "000000";
                          when "001001100110" => rgb <= "000000";
                          when "001001100111" => rgb <= "000000";
                          when "001001101000" => rgb <= "000000";
                          when "001001101001" => rgb <= "000000";
                          when "001010000000" => rgb <= "000000";
                          when "001010000001" => rgb <= "000000";
                          when "001010000010" => rgb <= "000000";
                          when "001010000011" => rgb <= "000000";
                          when "001010000100" => rgb <= "000000";
                          when "001010000101" => rgb <= "101000";
                          when "001010000110" => rgb <= "101000";
                          when "001010000111" => rgb <= "101000";
                          when "001010001000" => rgb <= "101000";
                          when "001010001001" => rgb <= "101000";
                          when "001010001010" => rgb <= "101000";
                          when "001010001011" => rgb <= "101000";
                          when "001010001100" => rgb <= "101000";
                          when "001010001101" => rgb <= "101000";
                          when "001010001110" => rgb <= "101000";
                          when "001010001111" => rgb <= "101000";
                          when "001010010000" => rgb <= "101000";
                          when "001010010001" => rgb <= "101000";
                          when "001010010010" => rgb <= "101000";
                          when "001010010011" => rgb <= "010000";
                          when "001010010100" => rgb <= "010000";
                          when "001010010101" => rgb <= "010000";
                          when "001010010110" => rgb <= "010000";
                          when "001010010111" => rgb <= "101000";
                          when "001010011000" => rgb <= "101000";
                          when "001010011001" => rgb <= "101000";
                          when "001010011010" => rgb <= "101000";
                          when "001010011011" => rgb <= "101000";
                          when "001010011100" => rgb <= "101000";
                          when "001010011101" => rgb <= "101000";
                          when "001010011110" => rgb <= "101000";
                          when "001010011111" => rgb <= "101000";
                          when "001010100000" => rgb <= "101000";
                          when "001010100001" => rgb <= "101000";
                          when "001010100010" => rgb <= "101000";
                          when "001010100011" => rgb <= "101000";
                          when "001010100100" => rgb <= "101000";
                          when "001010100101" => rgb <= "000000";
                          when "001010100110" => rgb <= "000000";
                          when "001010100111" => rgb <= "000000";
                          when "001010101000" => rgb <= "000000";
                          when "001010101001" => rgb <= "000000";
                          when "001011000000" => rgb <= "000000";
                          when "001011000001" => rgb <= "000000";
                          when "001011000010" => rgb <= "000000";
                          when "001011000011" => rgb <= "000000";
                          when "001011000100" => rgb <= "000000";
                          when "001011000101" => rgb <= "101000";
                          when "001011000110" => rgb <= "101000";
                          when "001011000111" => rgb <= "101000";
                          when "001011001000" => rgb <= "101000";
                          when "001011001001" => rgb <= "101000";
                          when "001011001010" => rgb <= "101000";
                          when "001011001011" => rgb <= "101000";
                          when "001011001100" => rgb <= "101000";
                          when "001011001101" => rgb <= "101000";
                          when "001011001110" => rgb <= "101000";
                          when "001011001111" => rgb <= "101000";
                          when "001011010000" => rgb <= "101000";
                          when "001011010001" => rgb <= "101000";
                          when "001011010010" => rgb <= "101000";
                          when "001011010011" => rgb <= "010000";
                          when "001011010100" => rgb <= "010000";
                          when "001011010101" => rgb <= "010000";
                          when "001011010110" => rgb <= "010000";
                          when "001011010111" => rgb <= "101000";
                          when "001011011000" => rgb <= "101000";
                          when "001011011001" => rgb <= "101000";
                          when "001011011010" => rgb <= "101000";
                          when "001011011011" => rgb <= "101000";
                          when "001011011100" => rgb <= "101000";
                          when "001011011101" => rgb <= "101000";
                          when "001011011110" => rgb <= "101000";
                          when "001011011111" => rgb <= "101000";
                          when "001011100000" => rgb <= "101000";
                          when "001011100001" => rgb <= "101000";
                          when "001011100010" => rgb <= "101000";
                          when "001011100011" => rgb <= "101000";
                          when "001011100100" => rgb <= "101000";
                          when "001011100101" => rgb <= "000000";
                          when "001011100110" => rgb <= "000000";
                          when "001011100111" => rgb <= "000000";
                          when "001011101000" => rgb <= "000000";
                          when "001011101001" => rgb <= "000000";
                          when "001100000000" => rgb <= "000000";
                          when "001100000001" => rgb <= "000000";
                          when "001100000010" => rgb <= "000000";
                          when "001100000011" => rgb <= "101000";
                          when "001100000100" => rgb <= "101000";
                          when "001100000101" => rgb <= "101000";
                          when "001100000110" => rgb <= "101000";
                          when "001100000111" => rgb <= "101000";
                          when "001100001000" => rgb <= "101001";
                          when "001100001001" => rgb <= "101001";
                          when "001100001010" => rgb <= "101001";
                          when "001100001011" => rgb <= "101001";
                          when "001100001100" => rgb <= "101001";
                          when "001100001101" => rgb <= "101001";
                          when "001100001110" => rgb <= "101000";
                          when "001100001111" => rgb <= "101000";
                          when "001100010000" => rgb <= "101000";
                          when "001100010001" => rgb <= "101000";
                          when "001100010010" => rgb <= "101000";
                          when "001100010011" => rgb <= "010000";
                          when "001100010100" => rgb <= "010000";
                          when "001100010101" => rgb <= "010000";
                          when "001100010110" => rgb <= "010000";
                          when "001100010111" => rgb <= "101000";
                          when "001100011000" => rgb <= "101000";
                          when "001100011001" => rgb <= "101000";
                          when "001100011010" => rgb <= "101000";
                          when "001100011011" => rgb <= "101000";
                          when "001100011100" => rgb <= "101000";
                          when "001100011101" => rgb <= "101000";
                          when "001100011110" => rgb <= "101000";
                          when "001100011111" => rgb <= "101000";
                          when "001100100000" => rgb <= "101000";
                          when "001100100001" => rgb <= "101000";
                          when "001100100010" => rgb <= "101000";
                          when "001100100011" => rgb <= "101000";
                          when "001100100100" => rgb <= "101000";
                          when "001100100101" => rgb <= "101000";
                          when "001100100110" => rgb <= "101000";
                          when "001100100111" => rgb <= "000000";
                          when "001100101000" => rgb <= "000000";
                          when "001100101001" => rgb <= "000000";
                          when "001101000000" => rgb <= "000000";
                          when "001101000001" => rgb <= "000000";
                          when "001101000010" => rgb <= "000000";
                          when "001101000011" => rgb <= "101000";
                          when "001101000100" => rgb <= "101000";
                          when "001101000101" => rgb <= "101000";
                          when "001101000110" => rgb <= "101000";
                          when "001101000111" => rgb <= "101000";
                          when "001101001000" => rgb <= "101001";
                          when "001101001001" => rgb <= "101001";
                          when "001101001010" => rgb <= "101001";
                          when "001101001011" => rgb <= "101001";
                          when "001101001100" => rgb <= "101001";
                          when "001101001101" => rgb <= "101001";
                          when "001101001110" => rgb <= "101000";
                          when "001101001111" => rgb <= "101000";
                          when "001101010000" => rgb <= "101000";
                          when "001101010001" => rgb <= "101000";
                          when "001101010010" => rgb <= "101000";
                          when "001101010011" => rgb <= "010000";
                          when "001101010100" => rgb <= "010000";
                          when "001101010101" => rgb <= "010000";
                          when "001101010110" => rgb <= "010000";
                          when "001101010111" => rgb <= "101000";
                          when "001101011000" => rgb <= "101000";
                          when "001101011001" => rgb <= "101000";
                          when "001101011010" => rgb <= "101000";
                          when "001101011011" => rgb <= "101000";
                          when "001101011100" => rgb <= "101000";
                          when "001101011101" => rgb <= "101000";
                          when "001101011110" => rgb <= "101000";
                          when "001101011111" => rgb <= "101000";
                          when "001101100000" => rgb <= "101000";
                          when "001101100001" => rgb <= "101000";
                          when "001101100010" => rgb <= "101000";
                          when "001101100011" => rgb <= "101000";
                          when "001101100100" => rgb <= "101000";
                          when "001101100101" => rgb <= "101000";
                          when "001101100110" => rgb <= "101000";
                          when "001101100111" => rgb <= "000000";
                          when "001101101000" => rgb <= "000000";
                          when "001101101001" => rgb <= "000000";
                          when "001110000000" => rgb <= "000000";
                          when "001110000001" => rgb <= "101001";
                          when "001110000010" => rgb <= "101000";
                          when "001110000011" => rgb <= "101000";
                          when "001110000100" => rgb <= "101000";
                          when "001110000101" => rgb <= "101000";
                          when "001110000110" => rgb <= "101000";
                          when "001110000111" => rgb <= "101001";
                          when "001110001000" => rgb <= "101001";
                          when "001110001001" => rgb <= "101001";
                          when "001110001010" => rgb <= "101000";
                          when "001110001011" => rgb <= "101000";
                          when "001110001100" => rgb <= "101000";
                          when "001110001101" => rgb <= "101000";
                          when "001110001110" => rgb <= "101000";
                          when "001110001111" => rgb <= "101000";
                          when "001110010000" => rgb <= "101000";
                          when "001110010001" => rgb <= "101000";
                          when "001110010010" => rgb <= "101000";
                          when "001110010011" => rgb <= "101000";
                          when "001110010100" => rgb <= "101000";
                          when "001110010101" => rgb <= "101000";
                          when "001110010110" => rgb <= "101000";
                          when "001110010111" => rgb <= "101000";
                          when "001110011000" => rgb <= "101000";
                          when "001110011001" => rgb <= "101000";
                          when "001110011010" => rgb <= "101000";
                          when "001110011011" => rgb <= "101000";
                          when "001110011100" => rgb <= "101000";
                          when "001110011101" => rgb <= "101000";
                          when "001110011110" => rgb <= "101000";
                          when "001110011111" => rgb <= "101000";
                          when "001110100000" => rgb <= "101000";
                          when "001110100001" => rgb <= "101000";
                          when "001110100010" => rgb <= "101000";
                          when "001110100011" => rgb <= "101000";
                          when "001110100100" => rgb <= "101000";
                          when "001110100101" => rgb <= "101000";
                          when "001110100110" => rgb <= "101000";
                          when "001110100111" => rgb <= "101000";
                          when "001110101000" => rgb <= "101001";
                          when "001110101001" => rgb <= "000000";
                          when "001111000000" => rgb <= "000000";
                          when "001111000001" => rgb <= "101001";
                          when "001111000010" => rgb <= "101000";
                          when "001111000011" => rgb <= "101000";
                          when "001111000100" => rgb <= "101000";
                          when "001111000101" => rgb <= "101001";
                          when "001111000110" => rgb <= "101001";
                          when "001111000111" => rgb <= "101001";
                          when "001111001000" => rgb <= "101001";
                          when "001111001001" => rgb <= "101001";
                          when "001111001010" => rgb <= "101000";
                          when "001111001011" => rgb <= "101000";
                          when "001111001100" => rgb <= "101000";
                          when "001111001101" => rgb <= "101000";
                          when "001111001110" => rgb <= "101000";
                          when "001111001111" => rgb <= "101000";
                          when "001111010000" => rgb <= "101000";
                          when "001111010001" => rgb <= "101000";
                          when "001111010010" => rgb <= "101000";
                          when "001111010011" => rgb <= "101000";
                          when "001111010100" => rgb <= "101000";
                          when "001111010101" => rgb <= "101000";
                          when "001111010110" => rgb <= "101000";
                          when "001111010111" => rgb <= "101000";
                          when "001111011000" => rgb <= "101000";
                          when "001111011001" => rgb <= "101000";
                          when "001111011010" => rgb <= "101000";
                          when "001111011011" => rgb <= "101000";
                          when "001111011100" => rgb <= "101000";
                          when "001111011101" => rgb <= "101000";
                          when "001111011110" => rgb <= "101000";
                          when "001111011111" => rgb <= "101000";
                          when "001111100000" => rgb <= "101000";
                          when "001111100001" => rgb <= "101000";
                          when "001111100010" => rgb <= "101000";
                          when "001111100011" => rgb <= "101000";
                          when "001111100100" => rgb <= "101000";
                          when "001111100101" => rgb <= "101000";
                          when "001111100110" => rgb <= "101000";
                          when "001111100111" => rgb <= "101000";
                          when "001111101000" => rgb <= "101000";
                          when "001111101001" => rgb <= "000000";
                          when "010000000000" => rgb <= "000000";
                          when "010000000001" => rgb <= "101001";
                          when "010000000010" => rgb <= "101000";
                          when "010000000011" => rgb <= "101000";
                          when "010000000100" => rgb <= "101000";
                          when "010000000101" => rgb <= "101001";
                          when "010000000110" => rgb <= "101001";
                          when "010000000111" => rgb <= "101001";
                          when "010000001000" => rgb <= "101001";
                          when "010000001001" => rgb <= "101000";
                          when "010000001010" => rgb <= "101000";
                          when "010000001011" => rgb <= "101000";
                          when "010000001100" => rgb <= "101000";
                          when "010000001101" => rgb <= "101000";
                          when "010000001110" => rgb <= "101000";
                          when "010000001111" => rgb <= "101000";
                          when "010000010000" => rgb <= "101000";
                          when "010000010001" => rgb <= "101000";
                          when "010000010010" => rgb <= "101000";
                          when "010000010011" => rgb <= "101000";
                          when "010000010100" => rgb <= "101000";
                          when "010000010101" => rgb <= "101000";
                          when "010000010110" => rgb <= "101000";
                          when "010000010111" => rgb <= "101000";
                          when "010000011000" => rgb <= "101000";
                          when "010000011001" => rgb <= "101000";
                          when "010000011010" => rgb <= "101000";
                          when "010000011011" => rgb <= "101000";
                          when "010000011100" => rgb <= "101000";
                          when "010000011101" => rgb <= "101000";
                          when "010000011110" => rgb <= "101000";
                          when "010000011111" => rgb <= "101000";
                          when "010000100000" => rgb <= "101000";
                          when "010000100001" => rgb <= "101000";
                          when "010000100010" => rgb <= "101000";
                          when "010000100011" => rgb <= "101000";
                          when "010000100100" => rgb <= "101000";
                          when "010000100101" => rgb <= "101000";
                          when "010000100110" => rgb <= "101000";
                          when "010000100111" => rgb <= "101000";
                          when "010000101000" => rgb <= "101000";
                          when "010000101001" => rgb <= "000000";
                          when "010001000000" => rgb <= "000000";
                          when "010001000001" => rgb <= "101001";
                          when "010001000010" => rgb <= "101000";
                          when "010001000011" => rgb <= "101000";
                          when "010001000100" => rgb <= "101000";
                          when "010001000101" => rgb <= "101001";
                          when "010001000110" => rgb <= "101001";
                          when "010001000111" => rgb <= "101001";
                          when "010001001000" => rgb <= "101000";
                          when "010001001001" => rgb <= "101000";
                          when "010001001010" => rgb <= "101000";
                          when "010001001011" => rgb <= "101000";
                          when "010001001100" => rgb <= "101000";
                          when "010001001101" => rgb <= "101000";
                          when "010001001110" => rgb <= "101000";
                          when "010001001111" => rgb <= "101000";
                          when "010001010000" => rgb <= "101000";
                          when "010001010001" => rgb <= "101000";
                          when "010001010010" => rgb <= "101000";
                          when "010001010011" => rgb <= "101000";
                          when "010001010100" => rgb <= "101000";
                          when "010001010101" => rgb <= "101000";
                          when "010001010110" => rgb <= "101000";
                          when "010001010111" => rgb <= "101000";
                          when "010001011000" => rgb <= "101000";
                          when "010001011001" => rgb <= "101000";
                          when "010001011010" => rgb <= "101000";
                          when "010001011011" => rgb <= "101000";
                          when "010001011100" => rgb <= "101000";
                          when "010001011101" => rgb <= "101000";
                          when "010001011110" => rgb <= "101000";
                          when "010001011111" => rgb <= "101000";
                          when "010001100000" => rgb <= "101000";
                          when "010001100001" => rgb <= "101000";
                          when "010001100010" => rgb <= "101000";
                          when "010001100011" => rgb <= "101000";
                          when "010001100100" => rgb <= "101000";
                          when "010001100101" => rgb <= "101000";
                          when "010001100110" => rgb <= "101000";
                          when "010001100111" => rgb <= "101000";
                          when "010001101000" => rgb <= "101001";
                          when "010001101001" => rgb <= "000000";
                          when "010010000000" => rgb <= "000000";
                          when "010010000001" => rgb <= "101001";
                          when "010010000010" => rgb <= "101000";
                          when "010010000011" => rgb <= "101000";
                          when "010010000100" => rgb <= "101000";
                          when "010010000101" => rgb <= "101001";
                          when "010010000110" => rgb <= "101001";
                          when "010010000111" => rgb <= "101000";
                          when "010010001000" => rgb <= "101000";
                          when "010010001001" => rgb <= "101000";
                          when "010010001010" => rgb <= "101000";
                          when "010010001011" => rgb <= "101000";
                          when "010010001100" => rgb <= "101000";
                          when "010010001101" => rgb <= "101000";
                          when "010010001110" => rgb <= "101000";
                          when "010010001111" => rgb <= "101000";
                          when "010010010000" => rgb <= "101000";
                          when "010010010001" => rgb <= "101000";
                          when "010010010010" => rgb <= "101000";
                          when "010010010011" => rgb <= "101000";
                          when "010010010100" => rgb <= "101000";
                          when "010010010101" => rgb <= "101000";
                          when "010010010110" => rgb <= "101000";
                          when "010010010111" => rgb <= "101000";
                          when "010010011000" => rgb <= "101000";
                          when "010010011001" => rgb <= "101000";
                          when "010010011010" => rgb <= "101000";
                          when "010010011011" => rgb <= "101000";
                          when "010010011100" => rgb <= "101000";
                          when "010010011101" => rgb <= "101000";
                          when "010010011110" => rgb <= "101000";
                          when "010010011111" => rgb <= "101000";
                          when "010010100000" => rgb <= "101000";
                          when "010010100001" => rgb <= "101000";
                          when "010010100010" => rgb <= "101000";
                          when "010010100011" => rgb <= "101000";
                          when "010010100100" => rgb <= "101000";
                          when "010010100101" => rgb <= "101000";
                          when "010010100110" => rgb <= "101000";
                          when "010010100111" => rgb <= "101000";
                          when "010010101000" => rgb <= "101000";
                          when "010010101001" => rgb <= "000000";
                          when "010011000000" => rgb <= "000000";
                          when "010011000001" => rgb <= "101001";
                          when "010011000010" => rgb <= "101000";
                          when "010011000011" => rgb <= "101000";
                          when "010011000100" => rgb <= "101000";
                          when "010011000101" => rgb <= "101001";
                          when "010011000110" => rgb <= "101001";
                          when "010011000111" => rgb <= "101000";
                          when "010011001000" => rgb <= "101000";
                          when "010011001001" => rgb <= "101000";
                          when "010011001010" => rgb <= "101000";
                          when "010011001011" => rgb <= "101000";
                          when "010011001100" => rgb <= "101000";
                          when "010011001101" => rgb <= "101000";
                          when "010011001110" => rgb <= "101000";
                          when "010011001111" => rgb <= "101000";
                          when "010011010000" => rgb <= "101000";
                          when "010011010001" => rgb <= "101000";
                          when "010011010010" => rgb <= "101000";
                          when "010011010011" => rgb <= "101000";
                          when "010011010100" => rgb <= "101000";
                          when "010011010101" => rgb <= "101000";
                          when "010011010110" => rgb <= "101000";
                          when "010011010111" => rgb <= "101000";
                          when "010011011000" => rgb <= "101000";
                          when "010011011001" => rgb <= "101000";
                          when "010011011010" => rgb <= "101000";
                          when "010011011011" => rgb <= "101000";
                          when "010011011100" => rgb <= "101000";
                          when "010011011101" => rgb <= "101000";
                          when "010011011110" => rgb <= "101000";
                          when "010011011111" => rgb <= "101000";
                          when "010011100000" => rgb <= "101000";
                          when "010011100001" => rgb <= "101000";
                          when "010011100010" => rgb <= "101000";
                          when "010011100011" => rgb <= "101000";
                          when "010011100100" => rgb <= "101000";
                          when "010011100101" => rgb <= "101000";
                          when "010011100110" => rgb <= "101000";
                          when "010011100111" => rgb <= "101000";
                          when "010011101000" => rgb <= "101000";
                          when "010011101001" => rgb <= "000000";
                          when "010100000000" => rgb <= "000000";
                          when "010100000001" => rgb <= "101001";
                          when "010100000010" => rgb <= "101000";
                          when "010100000011" => rgb <= "101000";
                          when "010100000100" => rgb <= "101000";
                          when "010100000101" => rgb <= "101001";
                          when "010100000110" => rgb <= "101001";
                          when "010100000111" => rgb <= "101000";
                          when "010100001000" => rgb <= "101000";
                          when "010100001001" => rgb <= "101000";
                          when "010100001010" => rgb <= "101000";
                          when "010100001011" => rgb <= "101000";
                          when "010100001100" => rgb <= "101000";
                          when "010100001101" => rgb <= "101000";
                          when "010100001110" => rgb <= "101000";
                          when "010100001111" => rgb <= "101000";
                          when "010100010000" => rgb <= "101000";
                          when "010100010001" => rgb <= "101000";
                          when "010100010010" => rgb <= "101000";
                          when "010100010011" => rgb <= "101000";
                          when "010100010100" => rgb <= "101000";
                          when "010100010101" => rgb <= "101000";
                          when "010100010110" => rgb <= "101000";
                          when "010100010111" => rgb <= "101000";
                          when "010100011000" => rgb <= "101000";
                          when "010100011001" => rgb <= "101000";
                          when "010100011010" => rgb <= "101000";
                          when "010100011011" => rgb <= "101000";
                          when "010100011100" => rgb <= "101000";
                          when "010100011101" => rgb <= "101000";
                          when "010100011110" => rgb <= "101000";
                          when "010100011111" => rgb <= "101000";
                          when "010100100000" => rgb <= "101000";
                          when "010100100001" => rgb <= "101000";
                          when "010100100010" => rgb <= "101000";
                          when "010100100011" => rgb <= "101000";
                          when "010100100100" => rgb <= "101000";
                          when "010100100101" => rgb <= "101000";
                          when "010100100110" => rgb <= "101000";
                          when "010100100111" => rgb <= "101000";
                          when "010100101000" => rgb <= "101000";
                          when "010100101001" => rgb <= "000000";
                          when "010101000000" => rgb <= "000000";
                          when "010101000001" => rgb <= "101001";
                          when "010101000010" => rgb <= "101000";
                          when "010101000011" => rgb <= "101000";
                          when "010101000100" => rgb <= "101000";
                          when "010101000101" => rgb <= "101000";
                          when "010101000110" => rgb <= "101000";
                          when "010101000111" => rgb <= "101000";
                          when "010101001000" => rgb <= "101000";
                          when "010101001001" => rgb <= "101000";
                          when "010101001010" => rgb <= "101000";
                          when "010101001011" => rgb <= "101000";
                          when "010101001100" => rgb <= "101000";
                          when "010101001101" => rgb <= "101000";
                          when "010101001110" => rgb <= "101000";
                          when "010101001111" => rgb <= "101000";
                          when "010101010000" => rgb <= "101000";
                          when "010101010001" => rgb <= "101000";
                          when "010101010010" => rgb <= "101000";
                          when "010101010011" => rgb <= "101000";
                          when "010101010100" => rgb <= "101000";
                          when "010101010101" => rgb <= "101000";
                          when "010101010110" => rgb <= "101000";
                          when "010101010111" => rgb <= "101000";
                          when "010101011000" => rgb <= "101000";
                          when "010101011001" => rgb <= "101000";
                          when "010101011010" => rgb <= "101000";
                          when "010101011011" => rgb <= "101000";
                          when "010101011100" => rgb <= "101000";
                          when "010101011101" => rgb <= "101000";
                          when "010101011110" => rgb <= "101000";
                          when "010101011111" => rgb <= "101000";
                          when "010101100000" => rgb <= "101000";
                          when "010101100001" => rgb <= "101000";
                          when "010101100010" => rgb <= "101000";
                          when "010101100011" => rgb <= "101000";
                          when "010101100100" => rgb <= "101000";
                          when "010101100101" => rgb <= "101000";
                          when "010101100110" => rgb <= "101000";
                          when "010101100111" => rgb <= "101000";
                          when "010101101000" => rgb <= "101000";
                          when "010101101001" => rgb <= "000000";
                          when "010110000000" => rgb <= "000000";
                          when "010110000001" => rgb <= "101001";
                          when "010110000010" => rgb <= "101000";
                          when "010110000011" => rgb <= "101000";
                          when "010110000100" => rgb <= "101000";
                          when "010110000101" => rgb <= "101000";
                          when "010110000110" => rgb <= "101000";
                          when "010110000111" => rgb <= "101000";
                          when "010110001000" => rgb <= "101000";
                          when "010110001001" => rgb <= "101000";
                          when "010110001010" => rgb <= "101000";
                          when "010110001011" => rgb <= "101000";
                          when "010110001100" => rgb <= "101000";
                          when "010110001101" => rgb <= "101000";
                          when "010110001110" => rgb <= "101000";
                          when "010110001111" => rgb <= "101000";
                          when "010110010000" => rgb <= "101000";
                          when "010110010001" => rgb <= "101000";
                          when "010110010010" => rgb <= "101000";
                          when "010110010011" => rgb <= "101000";
                          when "010110010100" => rgb <= "101000";
                          when "010110010101" => rgb <= "101000";
                          when "010110010110" => rgb <= "101000";
                          when "010110010111" => rgb <= "101000";
                          when "010110011000" => rgb <= "101000";
                          when "010110011001" => rgb <= "101000";
                          when "010110011010" => rgb <= "101000";
                          when "010110011011" => rgb <= "101000";
                          when "010110011100" => rgb <= "101000";
                          when "010110011101" => rgb <= "101000";
                          when "010110011110" => rgb <= "101000";
                          when "010110011111" => rgb <= "101000";
                          when "010110100000" => rgb <= "101000";
                          when "010110100001" => rgb <= "101000";
                          when "010110100010" => rgb <= "101000";
                          when "010110100011" => rgb <= "101000";
                          when "010110100100" => rgb <= "101000";
                          when "010110100101" => rgb <= "101000";
                          when "010110100110" => rgb <= "101000";
                          when "010110100111" => rgb <= "101000";
                          when "010110101000" => rgb <= "101001";
                          when "010110101001" => rgb <= "000000";
                          when "010111000000" => rgb <= "000000";
                          when "010111000001" => rgb <= "101001";
                          when "010111000010" => rgb <= "101000";
                          when "010111000011" => rgb <= "101000";
                          when "010111000100" => rgb <= "101000";
                          when "010111000101" => rgb <= "101000";
                          when "010111000110" => rgb <= "101000";
                          when "010111000111" => rgb <= "101000";
                          when "010111001000" => rgb <= "101000";
                          when "010111001001" => rgb <= "101000";
                          when "010111001010" => rgb <= "101000";
                          when "010111001011" => rgb <= "101000";
                          when "010111001100" => rgb <= "101000";
                          when "010111001101" => rgb <= "101000";
                          when "010111001110" => rgb <= "101000";
                          when "010111001111" => rgb <= "101000";
                          when "010111010000" => rgb <= "101000";
                          when "010111010001" => rgb <= "101000";
                          when "010111010010" => rgb <= "101000";
                          when "010111010011" => rgb <= "101000";
                          when "010111010100" => rgb <= "101000";
                          when "010111010101" => rgb <= "101000";
                          when "010111010110" => rgb <= "101000";
                          when "010111010111" => rgb <= "101000";
                          when "010111011000" => rgb <= "101000";
                          when "010111011001" => rgb <= "101000";
                          when "010111011010" => rgb <= "101000";
                          when "010111011011" => rgb <= "101000";
                          when "010111011100" => rgb <= "101000";
                          when "010111011101" => rgb <= "101000";
                          when "010111011110" => rgb <= "101000";
                          when "010111011111" => rgb <= "101000";
                          when "010111100000" => rgb <= "101000";
                          when "010111100001" => rgb <= "101000";
                          when "010111100010" => rgb <= "101000";
                          when "010111100011" => rgb <= "101000";
                          when "010111100100" => rgb <= "101000";
                          when "010111100101" => rgb <= "101000";
                          when "010111100110" => rgb <= "101000";
                          when "010111100111" => rgb <= "101000";
                          when "010111101000" => rgb <= "101001";
                          when "010111101001" => rgb <= "000000";
                          when "011000000000" => rgb <= "000000";
                          when "011000000001" => rgb <= "101001";
                          when "011000000010" => rgb <= "101000";
                          when "011000000011" => rgb <= "101000";
                          when "011000000100" => rgb <= "101000";
                          when "011000000101" => rgb <= "101000";
                          when "011000000110" => rgb <= "101000";
                          when "011000000111" => rgb <= "101000";
                          when "011000001000" => rgb <= "101000";
                          when "011000001001" => rgb <= "101000";
                          when "011000001010" => rgb <= "101000";
                          when "011000001011" => rgb <= "101000";
                          when "011000001100" => rgb <= "101000";
                          when "011000001101" => rgb <= "101000";
                          when "011000001110" => rgb <= "101000";
                          when "011000001111" => rgb <= "101000";
                          when "011000010000" => rgb <= "101000";
                          when "011000010001" => rgb <= "101000";
                          when "011000010010" => rgb <= "101000";
                          when "011000010011" => rgb <= "101000";
                          when "011000010100" => rgb <= "101000";
                          when "011000010101" => rgb <= "101000";
                          when "011000010110" => rgb <= "101000";
                          when "011000010111" => rgb <= "101000";
                          when "011000011000" => rgb <= "101000";
                          when "011000011001" => rgb <= "101000";
                          when "011000011010" => rgb <= "101000";
                          when "011000011011" => rgb <= "101000";
                          when "011000011100" => rgb <= "101000";
                          when "011000011101" => rgb <= "101000";
                          when "011000011110" => rgb <= "101000";
                          when "011000011111" => rgb <= "101000";
                          when "011000100000" => rgb <= "101000";
                          when "011000100001" => rgb <= "101000";
                          when "011000100010" => rgb <= "101000";
                          when "011000100011" => rgb <= "101000";
                          when "011000100100" => rgb <= "101000";
                          when "011000100101" => rgb <= "101000";
                          when "011000100110" => rgb <= "101000";
                          when "011000100111" => rgb <= "101000";
                          when "011000101000" => rgb <= "101001";
                          when "011000101001" => rgb <= "000000";
                          when "011001000000" => rgb <= "000000";
                          when "011001000001" => rgb <= "101001";
                          when "011001000010" => rgb <= "101000";
                          when "011001000011" => rgb <= "101000";
                          when "011001000100" => rgb <= "101000";
                          when "011001000101" => rgb <= "101000";
                          when "011001000110" => rgb <= "101000";
                          when "011001000111" => rgb <= "101000";
                          when "011001001000" => rgb <= "101000";
                          when "011001001001" => rgb <= "101000";
                          when "011001001010" => rgb <= "101000";
                          when "011001001011" => rgb <= "101000";
                          when "011001001100" => rgb <= "101000";
                          when "011001001101" => rgb <= "101000";
                          when "011001001110" => rgb <= "101000";
                          when "011001001111" => rgb <= "101000";
                          when "011001010000" => rgb <= "101000";
                          when "011001010001" => rgb <= "101000";
                          when "011001010010" => rgb <= "101000";
                          when "011001010011" => rgb <= "101000";
                          when "011001010100" => rgb <= "101000";
                          when "011001010101" => rgb <= "101000";
                          when "011001010110" => rgb <= "101000";
                          when "011001010111" => rgb <= "101000";
                          when "011001011000" => rgb <= "101000";
                          when "011001011001" => rgb <= "101000";
                          when "011001011010" => rgb <= "101000";
                          when "011001011011" => rgb <= "101000";
                          when "011001011100" => rgb <= "101000";
                          when "011001011101" => rgb <= "101000";
                          when "011001011110" => rgb <= "101000";
                          when "011001011111" => rgb <= "101000";
                          when "011001100000" => rgb <= "101000";
                          when "011001100001" => rgb <= "101000";
                          when "011001100010" => rgb <= "101000";
                          when "011001100011" => rgb <= "101000";
                          when "011001100100" => rgb <= "101000";
                          when "011001100101" => rgb <= "101000";
                          when "011001100110" => rgb <= "101000";
                          when "011001100111" => rgb <= "101000";
                          when "011001101000" => rgb <= "101001";
                          when "011001101001" => rgb <= "000000";
                          when "011010000000" => rgb <= "000000";
                          when "011010000001" => rgb <= "101001";
                          when "011010000010" => rgb <= "101000";
                          when "011010000011" => rgb <= "101000";
                          when "011010000100" => rgb <= "101000";
                          when "011010000101" => rgb <= "101000";
                          when "011010000110" => rgb <= "101000";
                          when "011010000111" => rgb <= "101000";
                          when "011010001000" => rgb <= "101000";
                          when "011010001001" => rgb <= "101000";
                          when "011010001010" => rgb <= "101000";
                          when "011010001011" => rgb <= "101000";
                          when "011010001100" => rgb <= "101000";
                          when "011010001101" => rgb <= "101000";
                          when "011010001110" => rgb <= "101000";
                          when "011010001111" => rgb <= "101000";
                          when "011010010000" => rgb <= "101000";
                          when "011010010001" => rgb <= "101000";
                          when "011010010010" => rgb <= "101000";
                          when "011010010011" => rgb <= "101000";
                          when "011010010100" => rgb <= "101000";
                          when "011010010101" => rgb <= "101000";
                          when "011010010110" => rgb <= "101000";
                          when "011010010111" => rgb <= "101000";
                          when "011010011000" => rgb <= "101000";
                          when "011010011001" => rgb <= "101000";
                          when "011010011010" => rgb <= "101000";
                          when "011010011011" => rgb <= "101000";
                          when "011010011100" => rgb <= "101000";
                          when "011010011101" => rgb <= "101000";
                          when "011010011110" => rgb <= "101000";
                          when "011010011111" => rgb <= "101000";
                          when "011010100000" => rgb <= "101000";
                          when "011010100001" => rgb <= "101000";
                          when "011010100010" => rgb <= "101000";
                          when "011010100011" => rgb <= "101000";
                          when "011010100100" => rgb <= "101000";
                          when "011010100101" => rgb <= "101000";
                          when "011010100110" => rgb <= "101000";
                          when "011010100111" => rgb <= "101000";
                          when "011010101000" => rgb <= "101001";
                          when "011010101001" => rgb <= "000000";
                          when "011011000000" => rgb <= "000000";
                          when "011011000001" => rgb <= "101001";
                          when "011011000010" => rgb <= "101000";
                          when "011011000011" => rgb <= "101000";
                          when "011011000100" => rgb <= "101000";
                          when "011011000101" => rgb <= "101000";
                          when "011011000110" => rgb <= "101000";
                          when "011011000111" => rgb <= "101000";
                          when "011011001000" => rgb <= "101000";
                          when "011011001001" => rgb <= "101000";
                          when "011011001010" => rgb <= "101000";
                          when "011011001011" => rgb <= "101000";
                          when "011011001100" => rgb <= "101000";
                          when "011011001101" => rgb <= "101000";
                          when "011011001110" => rgb <= "101000";
                          when "011011001111" => rgb <= "101000";
                          when "011011010000" => rgb <= "101000";
                          when "011011010001" => rgb <= "101000";
                          when "011011010010" => rgb <= "101000";
                          when "011011010011" => rgb <= "101000";
                          when "011011010100" => rgb <= "101000";
                          when "011011010101" => rgb <= "101000";
                          when "011011010110" => rgb <= "101000";
                          when "011011010111" => rgb <= "101000";
                          when "011011011000" => rgb <= "101000";
                          when "011011011001" => rgb <= "101000";
                          when "011011011010" => rgb <= "101000";
                          when "011011011011" => rgb <= "101000";
                          when "011011011100" => rgb <= "101000";
                          when "011011011101" => rgb <= "101000";
                          when "011011011110" => rgb <= "101000";
                          when "011011011111" => rgb <= "101000";
                          when "011011100000" => rgb <= "101000";
                          when "011011100001" => rgb <= "101000";
                          when "011011100010" => rgb <= "101000";
                          when "011011100011" => rgb <= "101000";
                          when "011011100100" => rgb <= "101000";
                          when "011011100101" => rgb <= "101000";
                          when "011011100110" => rgb <= "101000";
                          when "011011100111" => rgb <= "101000";
                          when "011011101000" => rgb <= "101001";
                          when "011011101001" => rgb <= "000000";
                          when "011100000000" => rgb <= "000000";
                          when "011100000001" => rgb <= "101001";
                          when "011100000010" => rgb <= "101000";
                          when "011100000011" => rgb <= "101000";
                          when "011100000100" => rgb <= "101000";
                          when "011100000101" => rgb <= "101000";
                          when "011100000110" => rgb <= "101000";
                          when "011100000111" => rgb <= "101000";
                          when "011100001000" => rgb <= "101000";
                          when "011100001001" => rgb <= "101000";
                          when "011100001010" => rgb <= "101000";
                          when "011100001011" => rgb <= "101000";
                          when "011100001100" => rgb <= "101000";
                          when "011100001101" => rgb <= "101000";
                          when "011100001110" => rgb <= "101000";
                          when "011100001111" => rgb <= "101000";
                          when "011100010000" => rgb <= "101000";
                          when "011100010001" => rgb <= "101000";
                          when "011100010010" => rgb <= "101000";
                          when "011100010011" => rgb <= "101000";
                          when "011100010100" => rgb <= "101000";
                          when "011100010101" => rgb <= "101000";
                          when "011100010110" => rgb <= "101000";
                          when "011100010111" => rgb <= "101000";
                          when "011100011000" => rgb <= "101000";
                          when "011100011001" => rgb <= "101000";
                          when "011100011010" => rgb <= "101000";
                          when "011100011011" => rgb <= "101000";
                          when "011100011100" => rgb <= "101000";
                          when "011100011101" => rgb <= "101000";
                          when "011100011110" => rgb <= "101000";
                          when "011100011111" => rgb <= "101000";
                          when "011100100000" => rgb <= "101000";
                          when "011100100001" => rgb <= "101000";
                          when "011100100010" => rgb <= "101000";
                          when "011100100011" => rgb <= "101000";
                          when "011100100100" => rgb <= "101000";
                          when "011100100101" => rgb <= "101000";
                          when "011100100110" => rgb <= "101000";
                          when "011100100111" => rgb <= "101000";
                          when "011100101000" => rgb <= "101001";
                          when "011100101001" => rgb <= "000000";
                          when "011101000000" => rgb <= "000000";
                          when "011101000001" => rgb <= "101001";
                          when "011101000010" => rgb <= "101000";
                          when "011101000011" => rgb <= "101000";
                          when "011101000100" => rgb <= "101000";
                          when "011101000101" => rgb <= "101000";
                          when "011101000110" => rgb <= "101000";
                          when "011101000111" => rgb <= "101000";
                          when "011101001000" => rgb <= "101000";
                          when "011101001001" => rgb <= "101000";
                          when "011101001010" => rgb <= "101000";
                          when "011101001011" => rgb <= "101000";
                          when "011101001100" => rgb <= "101000";
                          when "011101001101" => rgb <= "101000";
                          when "011101001110" => rgb <= "101000";
                          when "011101001111" => rgb <= "101000";
                          when "011101010000" => rgb <= "101000";
                          when "011101010001" => rgb <= "101000";
                          when "011101010010" => rgb <= "101000";
                          when "011101010011" => rgb <= "101000";
                          when "011101010100" => rgb <= "101000";
                          when "011101010101" => rgb <= "101000";
                          when "011101010110" => rgb <= "101000";
                          when "011101010111" => rgb <= "101000";
                          when "011101011000" => rgb <= "101000";
                          when "011101011001" => rgb <= "101000";
                          when "011101011010" => rgb <= "101000";
                          when "011101011011" => rgb <= "101000";
                          when "011101011100" => rgb <= "101000";
                          when "011101011101" => rgb <= "101000";
                          when "011101011110" => rgb <= "101000";
                          when "011101011111" => rgb <= "101000";
                          when "011101100000" => rgb <= "101000";
                          when "011101100001" => rgb <= "101000";
                          when "011101100010" => rgb <= "101000";
                          when "011101100011" => rgb <= "101000";
                          when "011101100100" => rgb <= "101000";
                          when "011101100101" => rgb <= "101000";
                          when "011101100110" => rgb <= "101000";
                          when "011101100111" => rgb <= "101000";
                          when "011101101000" => rgb <= "101001";
                          when "011101101001" => rgb <= "000000";
                          when "011110000000" => rgb <= "000000";
                          when "011110000001" => rgb <= "101001";
                          when "011110000010" => rgb <= "101000";
                          when "011110000011" => rgb <= "101000";
                          when "011110000100" => rgb <= "101000";
                          when "011110000101" => rgb <= "101000";
                          when "011110000110" => rgb <= "101000";
                          when "011110000111" => rgb <= "101000";
                          when "011110001000" => rgb <= "101000";
                          when "011110001001" => rgb <= "101000";
                          when "011110001010" => rgb <= "101000";
                          when "011110001011" => rgb <= "101000";
                          when "011110001100" => rgb <= "101000";
                          when "011110001101" => rgb <= "101000";
                          when "011110001110" => rgb <= "101000";
                          when "011110001111" => rgb <= "101000";
                          when "011110010000" => rgb <= "101000";
                          when "011110010001" => rgb <= "101000";
                          when "011110010010" => rgb <= "101000";
                          when "011110010011" => rgb <= "101000";
                          when "011110010100" => rgb <= "101000";
                          when "011110010101" => rgb <= "101000";
                          when "011110010110" => rgb <= "101000";
                          when "011110010111" => rgb <= "101000";
                          when "011110011000" => rgb <= "101000";
                          when "011110011001" => rgb <= "101000";
                          when "011110011010" => rgb <= "101000";
                          when "011110011011" => rgb <= "101000";
                          when "011110011100" => rgb <= "101000";
                          when "011110011101" => rgb <= "101000";
                          when "011110011110" => rgb <= "101000";
                          when "011110011111" => rgb <= "101000";
                          when "011110100000" => rgb <= "101000";
                          when "011110100001" => rgb <= "101000";
                          when "011110100010" => rgb <= "101000";
                          when "011110100011" => rgb <= "101000";
                          when "011110100100" => rgb <= "101000";
                          when "011110100101" => rgb <= "101000";
                          when "011110100110" => rgb <= "101000";
                          when "011110100111" => rgb <= "101000";
                          when "011110101000" => rgb <= "101001";
                          when "011110101001" => rgb <= "000000";
                          when "011111000000" => rgb <= "000000";
                          when "011111000001" => rgb <= "101001";
                          when "011111000010" => rgb <= "101000";
                          when "011111000011" => rgb <= "101000";
                          when "011111000100" => rgb <= "101000";
                          when "011111000101" => rgb <= "101000";
                          when "011111000110" => rgb <= "101000";
                          when "011111000111" => rgb <= "101000";
                          when "011111001000" => rgb <= "101000";
                          when "011111001001" => rgb <= "101000";
                          when "011111001010" => rgb <= "101000";
                          when "011111001011" => rgb <= "101000";
                          when "011111001100" => rgb <= "101000";
                          when "011111001101" => rgb <= "101000";
                          when "011111001110" => rgb <= "101000";
                          when "011111001111" => rgb <= "101000";
                          when "011111010000" => rgb <= "101000";
                          when "011111010001" => rgb <= "101000";
                          when "011111010010" => rgb <= "101000";
                          when "011111010011" => rgb <= "101000";
                          when "011111010100" => rgb <= "101000";
                          when "011111010101" => rgb <= "101000";
                          when "011111010110" => rgb <= "101000";
                          when "011111010111" => rgb <= "101000";
                          when "011111011000" => rgb <= "101000";
                          when "011111011001" => rgb <= "101000";
                          when "011111011010" => rgb <= "101000";
                          when "011111011011" => rgb <= "101000";
                          when "011111011100" => rgb <= "101000";
                          when "011111011101" => rgb <= "101000";
                          when "011111011110" => rgb <= "101000";
                          when "011111011111" => rgb <= "101000";
                          when "011111100000" => rgb <= "101000";
                          when "011111100001" => rgb <= "101000";
                          when "011111100010" => rgb <= "101000";
                          when "011111100011" => rgb <= "101000";
                          when "011111100100" => rgb <= "101000";
                          when "011111100101" => rgb <= "101000";
                          when "011111100110" => rgb <= "101000";
                          when "011111100111" => rgb <= "101000";
                          when "011111101000" => rgb <= "101001";
                          when "011111101001" => rgb <= "000000";
                          when "100000000000" => rgb <= "000000";
                          when "100000000001" => rgb <= "000000";
                          when "100000000010" => rgb <= "000000";
                          when "100000000011" => rgb <= "101000";
                          when "100000000100" => rgb <= "101000";
                          when "100000000101" => rgb <= "101000";
                          when "100000000110" => rgb <= "101000";
                          when "100000000111" => rgb <= "101000";
                          when "100000001000" => rgb <= "101000";
                          when "100000001001" => rgb <= "101000";
                          when "100000001010" => rgb <= "101000";
                          when "100000001011" => rgb <= "101000";
                          when "100000001100" => rgb <= "101000";
                          when "100000001101" => rgb <= "101000";
                          when "100000001110" => rgb <= "101000";
                          when "100000001111" => rgb <= "101000";
                          when "100000010000" => rgb <= "101000";
                          when "100000010001" => rgb <= "101000";
                          when "100000010010" => rgb <= "101000";
                          when "100000010011" => rgb <= "101000";
                          when "100000010100" => rgb <= "101000";
                          when "100000010101" => rgb <= "101000";
                          when "100000010110" => rgb <= "101000";
                          when "100000010111" => rgb <= "101000";
                          when "100000011000" => rgb <= "101000";
                          when "100000011001" => rgb <= "101000";
                          when "100000011010" => rgb <= "101000";
                          when "100000011011" => rgb <= "101000";
                          when "100000011100" => rgb <= "101000";
                          when "100000011101" => rgb <= "101000";
                          when "100000011110" => rgb <= "101000";
                          when "100000011111" => rgb <= "101000";
                          when "100000100000" => rgb <= "101000";
                          when "100000100001" => rgb <= "101000";
                          when "100000100010" => rgb <= "101000";
                          when "100000100011" => rgb <= "101000";
                          when "100000100100" => rgb <= "101000";
                          when "100000100101" => rgb <= "101000";
                          when "100000100110" => rgb <= "101000";
                          when "100000100111" => rgb <= "000000";
                          when "100000101000" => rgb <= "000000";
                          when "100000101001" => rgb <= "000000";
                          when "100001000000" => rgb <= "000000";
                          when "100001000001" => rgb <= "000000";
                          when "100001000010" => rgb <= "000000";
                          when "100001000011" => rgb <= "101000";
                          when "100001000100" => rgb <= "101000";
                          when "100001000101" => rgb <= "101000";
                          when "100001000110" => rgb <= "101000";
                          when "100001000111" => rgb <= "101000";
                          when "100001001000" => rgb <= "101000";
                          when "100001001001" => rgb <= "101000";
                          when "100001001010" => rgb <= "101000";
                          when "100001001011" => rgb <= "101000";
                          when "100001001100" => rgb <= "101000";
                          when "100001001101" => rgb <= "101000";
                          when "100001001110" => rgb <= "101000";
                          when "100001001111" => rgb <= "101000";
                          when "100001010000" => rgb <= "101000";
                          when "100001010001" => rgb <= "101000";
                          when "100001010010" => rgb <= "101000";
                          when "100001010011" => rgb <= "101000";
                          when "100001010100" => rgb <= "101000";
                          when "100001010101" => rgb <= "101000";
                          when "100001010110" => rgb <= "101000";
                          when "100001010111" => rgb <= "101000";
                          when "100001011000" => rgb <= "101000";
                          when "100001011001" => rgb <= "101000";
                          when "100001011010" => rgb <= "101000";
                          when "100001011011" => rgb <= "101000";
                          when "100001011100" => rgb <= "101000";
                          when "100001011101" => rgb <= "101000";
                          when "100001011110" => rgb <= "101000";
                          when "100001011111" => rgb <= "101000";
                          when "100001100000" => rgb <= "101000";
                          when "100001100001" => rgb <= "101000";
                          when "100001100010" => rgb <= "101000";
                          when "100001100011" => rgb <= "101000";
                          when "100001100100" => rgb <= "101000";
                          when "100001100101" => rgb <= "101000";
                          when "100001100110" => rgb <= "101000";
                          when "100001100111" => rgb <= "000000";
                          when "100001101000" => rgb <= "000000";
                          when "100001101001" => rgb <= "000000";
                          when "100010000000" => rgb <= "000000";
                          when "100010000001" => rgb <= "000000";
                          when "100010000010" => rgb <= "000000";
                          when "100010000011" => rgb <= "101000";
                          when "100010000100" => rgb <= "101000";
                          when "100010000101" => rgb <= "101000";
                          when "100010000110" => rgb <= "101000";
                          when "100010000111" => rgb <= "101000";
                          when "100010001000" => rgb <= "101000";
                          when "100010001001" => rgb <= "101000";
                          when "100010001010" => rgb <= "101000";
                          when "100010001011" => rgb <= "101000";
                          when "100010001100" => rgb <= "101000";
                          when "100010001101" => rgb <= "101000";
                          when "100010001110" => rgb <= "101000";
                          when "100010001111" => rgb <= "101000";
                          when "100010010000" => rgb <= "101000";
                          when "100010010001" => rgb <= "101000";
                          when "100010010010" => rgb <= "101000";
                          when "100010010011" => rgb <= "101000";
                          when "100010010100" => rgb <= "101000";
                          when "100010010101" => rgb <= "101000";
                          when "100010010110" => rgb <= "101000";
                          when "100010010111" => rgb <= "101000";
                          when "100010011000" => rgb <= "101000";
                          when "100010011001" => rgb <= "101000";
                          when "100010011010" => rgb <= "101000";
                          when "100010011011" => rgb <= "101000";
                          when "100010011100" => rgb <= "101000";
                          when "100010011101" => rgb <= "101000";
                          when "100010011110" => rgb <= "101000";
                          when "100010011111" => rgb <= "101000";
                          when "100010100000" => rgb <= "101000";
                          when "100010100001" => rgb <= "101000";
                          when "100010100010" => rgb <= "101000";
                          when "100010100011" => rgb <= "101000";
                          when "100010100100" => rgb <= "101000";
                          when "100010100101" => rgb <= "101000";
                          when "100010100110" => rgb <= "101000";
                          when "100010100111" => rgb <= "000000";
                          when "100010101000" => rgb <= "000000";
                          when "100010101001" => rgb <= "000000";
                          when "100011000000" => rgb <= "000000";
                          when "100011000001" => rgb <= "000000";
                          when "100011000010" => rgb <= "000000";
                          when "100011000011" => rgb <= "101000";
                          when "100011000100" => rgb <= "101000";
                          when "100011000101" => rgb <= "101000";
                          when "100011000110" => rgb <= "101000";
                          when "100011000111" => rgb <= "101000";
                          when "100011001000" => rgb <= "101000";
                          when "100011001001" => rgb <= "101000";
                          when "100011001010" => rgb <= "101000";
                          when "100011001011" => rgb <= "101000";
                          when "100011001100" => rgb <= "101000";
                          when "100011001101" => rgb <= "101000";
                          when "100011001110" => rgb <= "101000";
                          when "100011001111" => rgb <= "101000";
                          when "100011010000" => rgb <= "101000";
                          when "100011010001" => rgb <= "101000";
                          when "100011010010" => rgb <= "101000";
                          when "100011010011" => rgb <= "101000";
                          when "100011010100" => rgb <= "101000";
                          when "100011010101" => rgb <= "101000";
                          when "100011010110" => rgb <= "101000";
                          when "100011010111" => rgb <= "101000";
                          when "100011011000" => rgb <= "101000";
                          when "100011011001" => rgb <= "101000";
                          when "100011011010" => rgb <= "101000";
                          when "100011011011" => rgb <= "101000";
                          when "100011011100" => rgb <= "101000";
                          when "100011011101" => rgb <= "101000";
                          when "100011011110" => rgb <= "101000";
                          when "100011011111" => rgb <= "101000";
                          when "100011100000" => rgb <= "101000";
                          when "100011100001" => rgb <= "101000";
                          when "100011100010" => rgb <= "101000";
                          when "100011100011" => rgb <= "101000";
                          when "100011100100" => rgb <= "101000";
                          when "100011100101" => rgb <= "101000";
                          when "100011100110" => rgb <= "101000";
                          when "100011100111" => rgb <= "000000";
                          when "100011101000" => rgb <= "000000";
                          when "100011101001" => rgb <= "000000";
                          when "100100000000" => rgb <= "000000";
                          when "100100000001" => rgb <= "000000";
                          when "100100000010" => rgb <= "000000";
                          when "100100000011" => rgb <= "000000";
                          when "100100000100" => rgb <= "000000";
                          when "100100000101" => rgb <= "101000";
                          when "100100000110" => rgb <= "101000";
                          when "100100000111" => rgb <= "101000";
                          when "100100001000" => rgb <= "101000";
                          when "100100001001" => rgb <= "101000";
                          when "100100001010" => rgb <= "101000";
                          when "100100001011" => rgb <= "101000";
                          when "100100001100" => rgb <= "101000";
                          when "100100001101" => rgb <= "101000";
                          when "100100001110" => rgb <= "101000";
                          when "100100001111" => rgb <= "101000";
                          when "100100010000" => rgb <= "101000";
                          when "100100010001" => rgb <= "101000";
                          when "100100010010" => rgb <= "101000";
                          when "100100010011" => rgb <= "101000";
                          when "100100010100" => rgb <= "101000";
                          when "100100010101" => rgb <= "101000";
                          when "100100010110" => rgb <= "101000";
                          when "100100010111" => rgb <= "101000";
                          when "100100011000" => rgb <= "101000";
                          when "100100011001" => rgb <= "101000";
                          when "100100011010" => rgb <= "101000";
                          when "100100011011" => rgb <= "101000";
                          when "100100011100" => rgb <= "101000";
                          when "100100011101" => rgb <= "101000";
                          when "100100011110" => rgb <= "101000";
                          when "100100011111" => rgb <= "101000";
                          when "100100100000" => rgb <= "101000";
                          when "100100100001" => rgb <= "101000";
                          when "100100100010" => rgb <= "101000";
                          when "100100100011" => rgb <= "101000";
                          when "100100100100" => rgb <= "101000";
                          when "100100100101" => rgb <= "000000";
                          when "100100100110" => rgb <= "000000";
                          when "100100100111" => rgb <= "000000";
                          when "100100101000" => rgb <= "000000";
                          when "100100101001" => rgb <= "000000";
                          when "100101000000" => rgb <= "000000";
                          when "100101000001" => rgb <= "000000";
                          when "100101000010" => rgb <= "000000";
                          when "100101000011" => rgb <= "000000";
                          when "100101000100" => rgb <= "000000";
                          when "100101000101" => rgb <= "000000";
                          when "100101000110" => rgb <= "101000";
                          when "100101000111" => rgb <= "101000";
                          when "100101001000" => rgb <= "101000";
                          when "100101001001" => rgb <= "101000";
                          when "100101001010" => rgb <= "101000";
                          when "100101001011" => rgb <= "101000";
                          when "100101001100" => rgb <= "101000";
                          when "100101001101" => rgb <= "101000";
                          when "100101001110" => rgb <= "101000";
                          when "100101001111" => rgb <= "101000";
                          when "100101010000" => rgb <= "101000";
                          when "100101010001" => rgb <= "101000";
                          when "100101010010" => rgb <= "101000";
                          when "100101010011" => rgb <= "101000";
                          when "100101010100" => rgb <= "101000";
                          when "100101010101" => rgb <= "101000";
                          when "100101010110" => rgb <= "101000";
                          when "100101010111" => rgb <= "101000";
                          when "100101011000" => rgb <= "101000";
                          when "100101011001" => rgb <= "101000";
                          when "100101011010" => rgb <= "101000";
                          when "100101011011" => rgb <= "101000";
                          when "100101011100" => rgb <= "101000";
                          when "100101011101" => rgb <= "101000";
                          when "100101011110" => rgb <= "101000";
                          when "100101011111" => rgb <= "101000";
                          when "100101100000" => rgb <= "101000";
                          when "100101100001" => rgb <= "101000";
                          when "100101100010" => rgb <= "101000";
                          when "100101100011" => rgb <= "101000";
                          when "100101100100" => rgb <= "000000";
                          when "100101100101" => rgb <= "000000";
                          when "100101100110" => rgb <= "000000";
                          when "100101100111" => rgb <= "000000";
                          when "100101101000" => rgb <= "000000";
                          when "100101101001" => rgb <= "000000";
                          when "100110000000" => rgb <= "000000";
                          when "100110000001" => rgb <= "000000";
                          when "100110000010" => rgb <= "000000";
                          when "100110000011" => rgb <= "000000";
                          when "100110000100" => rgb <= "000000";
                          when "100110000101" => rgb <= "000000";
                          when "100110000110" => rgb <= "101000";
                          when "100110000111" => rgb <= "101000";
                          when "100110001000" => rgb <= "101000";
                          when "100110001001" => rgb <= "101000";
                          when "100110001010" => rgb <= "101000";
                          when "100110001011" => rgb <= "101000";
                          when "100110001100" => rgb <= "101000";
                          when "100110001101" => rgb <= "101000";
                          when "100110001110" => rgb <= "101000";
                          when "100110001111" => rgb <= "101000";
                          when "100110010000" => rgb <= "101000";
                          when "100110010001" => rgb <= "101000";
                          when "100110010010" => rgb <= "101000";
                          when "100110010011" => rgb <= "101000";
                          when "100110010100" => rgb <= "101000";
                          when "100110010101" => rgb <= "101000";
                          when "100110010110" => rgb <= "101000";
                          when "100110010111" => rgb <= "101000";
                          when "100110011000" => rgb <= "101000";
                          when "100110011001" => rgb <= "101000";
                          when "100110011010" => rgb <= "101000";
                          when "100110011011" => rgb <= "101000";
                          when "100110011100" => rgb <= "101000";
                          when "100110011101" => rgb <= "101000";
                          when "100110011110" => rgb <= "101000";
                          when "100110011111" => rgb <= "101000";
                          when "100110100000" => rgb <= "101000";
                          when "100110100001" => rgb <= "101000";
                          when "100110100010" => rgb <= "101000";
                          when "100110100011" => rgb <= "101000";
                          when "100110100100" => rgb <= "000000";
                          when "100110100101" => rgb <= "000000";
                          when "100110100110" => rgb <= "000000";
                          when "100110100111" => rgb <= "000000";
                          when "100110101000" => rgb <= "000000";
                          when "100110101001" => rgb <= "000000";
                          when "100111000000" => rgb <= "000000";
                          when "100111000001" => rgb <= "000000";
                          when "100111000010" => rgb <= "000000";
                          when "100111000011" => rgb <= "000000";
                          when "100111000100" => rgb <= "000000";
                          when "100111000101" => rgb <= "000000";
                          when "100111000110" => rgb <= "000000";
                          when "100111000111" => rgb <= "000000";
                          when "100111001000" => rgb <= "000000";
                          when "100111001001" => rgb <= "000000";
                          when "100111001010" => rgb <= "101000";
                          when "100111001011" => rgb <= "101000";
                          when "100111001100" => rgb <= "101000";
                          when "100111001101" => rgb <= "101000";
                          when "100111001110" => rgb <= "101000";
                          when "100111001111" => rgb <= "101000";
                          when "100111010000" => rgb <= "101000";
                          when "100111010001" => rgb <= "101000";
                          when "100111010010" => rgb <= "101000";
                          when "100111010011" => rgb <= "000000";
                          when "100111010100" => rgb <= "000000";
                          when "100111010101" => rgb <= "000000";
                          when "100111010110" => rgb <= "000000";
                          when "100111010111" => rgb <= "101000";
                          when "100111011000" => rgb <= "101000";
                          when "100111011001" => rgb <= "101000";
                          when "100111011010" => rgb <= "101000";
                          when "100111011011" => rgb <= "101000";
                          when "100111011100" => rgb <= "101000";
                          when "100111011101" => rgb <= "101000";
                          when "100111011110" => rgb <= "101000";
                          when "100111011111" => rgb <= "101000";
                          when "100111100000" => rgb <= "000000";
                          when "100111100001" => rgb <= "000000";
                          when "100111100010" => rgb <= "000000";
                          when "100111100011" => rgb <= "000000";
                          when "100111100100" => rgb <= "000000";
                          when "100111100101" => rgb <= "000000";
                          when "100111100110" => rgb <= "000000";
                          when "100111100111" => rgb <= "000000";
                          when "100111101000" => rgb <= "000000";
                          when "100111101001" => rgb <= "000000";
                          when "101000000000" => rgb <= "000000";
                          when "101000000001" => rgb <= "000000";
                          when "101000000010" => rgb <= "000000";
                          when "101000000011" => rgb <= "000000";
                          when "101000000100" => rgb <= "000000";
                          when "101000000101" => rgb <= "000000";
                          when "101000000110" => rgb <= "000000";
                          when "101000000111" => rgb <= "000000";
                          when "101000001000" => rgb <= "000000";
                          when "101000001001" => rgb <= "000000";
                          when "101000001010" => rgb <= "101001";
                          when "101000001011" => rgb <= "101001";
                          when "101000001100" => rgb <= "101000";
                          when "101000001101" => rgb <= "101001";
                          when "101000001110" => rgb <= "101001";
                          when "101000001111" => rgb <= "101000";
                          when "101000010000" => rgb <= "101000";
                          when "101000010001" => rgb <= "101001";
                          when "101000010010" => rgb <= "101000";
                          when "101000010011" => rgb <= "000000";
                          when "101000010100" => rgb <= "000000";
                          when "101000010101" => rgb <= "000000";
                          when "101000010110" => rgb <= "000000";
                          when "101000010111" => rgb <= "101001";
                          when "101000011000" => rgb <= "101001";
                          when "101000011001" => rgb <= "101001";
                          when "101000011010" => rgb <= "101001";
                          when "101000011011" => rgb <= "101001";
                          when "101000011100" => rgb <= "101001";
                          when "101000011101" => rgb <= "101001";
                          when "101000011110" => rgb <= "101001";
                          when "101000011111" => rgb <= "101001";
                          when "101000100000" => rgb <= "000000";
                          when "101000100001" => rgb <= "000000";
                          when "101000100010" => rgb <= "000000";
                          when "101000100011" => rgb <= "000000";
                          when "101000100100" => rgb <= "000000";
                          when "101000100101" => rgb <= "000000";
                          when "101000100110" => rgb <= "000000";
                          when "101000100111" => rgb <= "000000";
                          when "101000101000" => rgb <= "000000";
                          when "101000101001" => rgb <= "000000";
                          when "101001000000" => rgb <= "000000";
                          when "101001000001" => rgb <= "000000";
                          when "101001000010" => rgb <= "000000";
                          when "101001000011" => rgb <= "000000";
                          when "101001000100" => rgb <= "000000";
                          when "101001000101" => rgb <= "000000";
                          when "101001000110" => rgb <= "000000";
                          when "101001000111" => rgb <= "000000";
                          when "101001001000" => rgb <= "000000";
                          when "101001001001" => rgb <= "000000";
                          when "101001001010" => rgb <= "000000";
                          when "101001001011" => rgb <= "000000";
                          when "101001001100" => rgb <= "000000";
                          when "101001001101" => rgb <= "000000";
                          when "101001001110" => rgb <= "000000";
                          when "101001001111" => rgb <= "000000";
                          when "101001010000" => rgb <= "000000";
                          when "101001010001" => rgb <= "000000";
                          when "101001010010" => rgb <= "000000";
                          when "101001010011" => rgb <= "000000";
                          when "101001010100" => rgb <= "000000";
                          when "101001010101" => rgb <= "000000";
                          when "101001010110" => rgb <= "000000";
                          when "101001010111" => rgb <= "000000";
                          when "101001011000" => rgb <= "000000";
                          when "101001011001" => rgb <= "000000";
                          when "101001011010" => rgb <= "000000";
                          when "101001011011" => rgb <= "000000";
                          when "101001011100" => rgb <= "000000";
                          when "101001011101" => rgb <= "000000";
                          when "101001011110" => rgb <= "000000";
                          when "101001011111" => rgb <= "000000";
                          when "101001100000" => rgb <= "000000";
                          when "101001100001" => rgb <= "000000";
                          when "101001100010" => rgb <= "000000";
                          when "101001100011" => rgb <= "000000";
                          when "101001100100" => rgb <= "000000";
                          when "101001100101" => rgb <= "000000";
                          when "101001100110" => rgb <= "000000";
                          when "101001100111" => rgb <= "000000";
                          when "101001101000" => rgb <= "000000";
                          when "101001101001" => rgb <= "000000";
                              when others => rgb <= "000000";
                end case;
				else
					rgb <= "000000";
				end if;
            end if;
            end process;
        end;
                
