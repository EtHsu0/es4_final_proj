library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity top is 
  port(
        -- NES controllers input
        -- VGA display output
  );
end top;

architecture synth of top is
-- Components for VGA
-- Components for NES?
-- Components for Snake
-- Components for menu selection?
-- Components for setting options
-- Components for random apples generation 
        -- (Maybe component will be called in another component)
        -- Return different combinations of settings.
        -- Bitpacking information into 
-- State we have? Initial state (Menu selection)
        -- One state for each menu options (Start, Settings, End)
        -- Other "sub" states for each options
                -- For example after start, we have ongoing, game over, etc.
begin
--     a <= '1';
end;



